#=============================================================================
# LEF - UNIT CELL
# Copyright (c) 2008 FUJITSU MICROELECTRONICS LIMITED  All rights reserved.
#=============================================================================
# LIBRARY        : CS202SN (CS202 9-track height cell) ;
# CLASSIFICATION : CUSTOM SET (LPDK) ;
# FILETYPE       : LEF ;
# DATE           : 2008/04/04 ;
# REVISION       : 1.1 ;
# DESIGNER       : A.NISHIWAKI (FUJITSU VLSI LIMITED) ;
# SOURCE         : cs202sn_uc_lpdk.gds_r01p1.gds ;
#
#=============================================================================
# HISTORY
#=============================================================================
# Rev.  Date(YMD)   Comment
# ----  ----------  ----------------------------------------------------------
# 1.1   2008/04/04  Official Release [ 24 cell ]
#                   [mod] 24 cells
#                   Add Well layer | Optimize Antenna parameter
# 1.0   2007/07/20  Official Release [ 24 cell ]
#                   [add] 24 cells

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

MACRO SC22AOBWSCLXL1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22AOBWSCLXL1 0 0 ;
  SIZE 4.6 BY 3.6 ;
  SYMMETRY X Y ;
  SITE WCORE3600 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.0735 LAYER MET1 ;
    ANTENNAMAXCUTCAR 40.819562 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDDG ;
    PORT
      LAYER MET1 ;
        RECT 1.635 0.4 1.735 0.85 ;
        RECT 1.635 0.75 2.435 0.85 ;
      LAYER CUT01 ;
        RECT 1.64 0.45 1.73 0.54 ;
        RECT 2.3 0.755 2.39 0.845 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 0.5 2.82 ;
        RECT 4.1 0.78 5.1 2.82 ;
      LAYER MET1 ;
        RECT 0 1.64 4.6 1.96 ;
      LAYER CUT01 ;
        RECT 0.175 1.86 0.265 1.95 ;
        RECT 0.175 1.65 0.265 1.74 ;
        RECT 4.335 1.86 4.425 1.95 ;
        RECT 4.335 1.65 4.425 1.74 ;
    END
  END VDD
  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT 1.5 0.78 3.1 2.82 ;
      LAYER MET1 ;
        RECT 1.8 2.125 1.9 2.46 ;
        RECT 2.32 2.125 2.42 2.46 ;
        RECT 2.84 2.125 2.94 2.46 ;
        RECT 0.06 2.125 4.54 2.275 ;
        RECT 1.675 1.14 1.775 1.475 ;
        RECT 2.02 1.12 2.12 1.475 ;
        RECT 0.06 1.325 4.54 1.475 ;
      LAYER CUT01 ;
        RECT 1.68 1.38 1.77 1.47 ;
        RECT 1.68 1.18 1.77 1.27 ;
        RECT 1.805 2.33 1.895 2.42 ;
        RECT 1.805 2.13 1.895 2.22 ;
        RECT 2.025 1.36 2.115 1.45 ;
        RECT 2.025 1.16 2.115 1.25 ;
        RECT 2.325 2.33 2.415 2.42 ;
        RECT 2.325 2.13 2.415 2.22 ;
        RECT 2.545 1.355 2.635 1.445 ;
        RECT 2.845 2.33 2.935 2.42 ;
        RECT 2.845 2.13 2.935 2.22 ;
    END
  END VDDG
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 2.32 3.04 2.42 3.76 ;
        RECT 2.84 3.04 2.94 3.76 ;
        RECT 0 3.44 4.6 3.76 ;
        RECT 2.28 -0.16 2.38 0.555 ;
        RECT 0 -0.16 4.6 0.16 ;
      LAYER CUT01 ;
        RECT 2.285 0.425 2.375 0.515 ;
        RECT 2.285 0.225 2.375 0.315 ;
        RECT 2.325 3.28 2.415 3.37 ;
        RECT 2.325 3.08 2.415 3.17 ;
        RECT 2.845 3.28 2.935 3.37 ;
        RECT 2.845 3.08 2.935 3.17 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4477 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 2.025 2.415 2.195 3.3 ;
        RECT 2.025 2.7 2.715 2.9 ;
        RECT 2.545 2.415 2.715 3.3 ;
      LAYER CUT01 ;
        RECT 2.065 3.205 2.155 3.295 ;
        RECT 2.065 3.005 2.155 3.095 ;
        RECT 2.065 2.455 2.155 2.545 ;
        RECT 2.585 3.205 2.675 3.295 ;
        RECT 2.585 3.005 2.675 3.095 ;
        RECT 2.585 2.455 2.675 2.545 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT 0.5 -0.5 1.5 4.1 ;
        RECT 3.1 -0.5 4.1 4.1 ;
        RECT -0.5 -0.5 5.1 0.78 ;
        RECT -0.5 2.82 5.1 4.1 ;
    END
  END VPW
  OBS
    LAYER MET1 ;
      RECT 2.54 0.29 2.64 1.205 ;
      RECT 2.24 1.105 2.875 1.205 ;
  END
END SC22AOBWSCLXL1

MACRO SC22AOBWSCLXP1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22AOBWSCLXP1 0 0 ;
  SIZE 5.2 BY 3.6 ;
  SYMMETRY X Y ;
  SITE WCORE3600 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.15375 LAYER MET1 ;
    ANTENNAMAXCUTCAR 39.027566 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDDG ;
    PORT
      LAYER MET1 ;
        RECT 1.635 0.4 1.735 0.85 ;
        RECT 1.635 0.73 2.715 0.85 ;
      LAYER CUT01 ;
        RECT 1.64 0.45 1.73 0.54 ;
        RECT 2.315 0.73 2.405 0.82 ;
        RECT 2.575 0.73 2.665 0.82 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 0.5 2.82 ;
        RECT 4.7 0.78 5.7 2.82 ;
      LAYER MET1 ;
        RECT 0 1.64 5.2 1.96 ;
      LAYER CUT01 ;
        RECT 0.175 1.86 0.265 1.95 ;
        RECT 0.175 1.65 0.265 1.74 ;
        RECT 4.935 1.86 5.025 1.95 ;
        RECT 4.935 1.65 5.025 1.74 ;
    END
  END VDD
  PIN VDDG
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT 1.5 0.78 3.7 2.82 ;
      LAYER MET1 ;
        RECT 1.79 2.125 1.89 2.46 ;
        RECT 3.42 2.125 3.52 2.46 ;
        RECT 0.06 2.125 5.14 2.275 ;
        RECT 1.675 1.14 1.775 1.475 ;
        RECT 3.42 1.14 3.52 1.475 ;
        RECT 0.06 1.325 5.14 1.475 ;
      LAYER CUT01 ;
        RECT 1.68 1.38 1.77 1.47 ;
        RECT 1.68 1.18 1.77 1.27 ;
        RECT 1.795 2.33 1.885 2.42 ;
        RECT 1.795 2.13 1.885 2.22 ;
        RECT 2.315 2.155 2.405 2.245 ;
        RECT 2.315 1.355 2.405 1.445 ;
        RECT 2.835 2.155 2.925 2.245 ;
        RECT 2.835 1.355 2.925 1.445 ;
        RECT 3.425 2.33 3.515 2.42 ;
        RECT 3.425 2.13 3.515 2.22 ;
        RECT 3.425 1.38 3.515 1.47 ;
        RECT 3.425 1.18 3.515 1.27 ;
    END
  END VDDG
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 1.79 3.03 1.89 3.76 ;
        RECT 2.31 3.03 2.41 3.76 ;
        RECT 2.83 3.03 2.93 3.76 ;
        RECT 3.42 3.03 3.52 3.76 ;
        RECT 0 3.44 5.2 3.76 ;
        RECT 2.31 -0.16 2.41 0.55 ;
        RECT 2.83 -0.16 2.93 0.38 ;
        RECT 0 -0.16 5.2 0.16 ;
      LAYER CUT01 ;
        RECT 1.795 3.28 1.885 3.37 ;
        RECT 1.795 3.07 1.885 3.16 ;
        RECT 2.315 3.28 2.405 3.37 ;
        RECT 2.315 3.07 2.405 3.16 ;
        RECT 2.315 0.42 2.405 0.51 ;
        RECT 2.315 0.21 2.405 0.3 ;
        RECT 2.835 3.28 2.925 3.37 ;
        RECT 2.835 3.07 2.925 3.16 ;
        RECT 2.835 0.24 2.925 0.33 ;
        RECT 3.425 3.28 3.515 3.37 ;
        RECT 3.425 3.07 3.515 3.16 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.0063 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 2.015 2.415 2.185 3.3 ;
        RECT 2.535 2.415 2.705 3.3 ;
        RECT 2.015 2.55 3.26 2.85 ;
        RECT 3.09 2.415 3.26 3.3 ;
      LAYER CUT01 ;
        RECT 2.055 3.205 2.145 3.295 ;
        RECT 2.055 3.005 2.145 3.095 ;
        RECT 2.055 2.455 2.145 2.545 ;
        RECT 2.575 3.205 2.665 3.295 ;
        RECT 2.575 3.005 2.665 3.095 ;
        RECT 2.575 2.455 2.665 2.545 ;
        RECT 3.13 3.205 3.22 3.295 ;
        RECT 3.13 3.005 3.22 3.095 ;
        RECT 3.13 2.455 3.22 2.545 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT 0.5 -0.5 1.5 4.1 ;
        RECT 3.7 -0.5 4.7 4.1 ;
        RECT -0.5 -0.5 5.7 0.78 ;
        RECT -0.5 2.82 5.7 4.1 ;
    END
  END VPW
  OBS
    LAYER MET1 ;
      RECT 2.57 0.285 2.67 0.62 ;
      RECT 2.53 0.52 3.11 0.62 ;
      RECT 3.01 0.715 3.485 0.815 ;
      RECT 3.01 0.52 3.11 1.15 ;
      RECT 2.005 1.05 3.11 1.15 ;
  END
END SC22AOBWSCLXP1

MACRO SC22ISOANDCLXL1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22ISOANDCLXL1 0 0 ;
  SIZE 2.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE CORE1800 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.117 LAYER MET1 ;
    ANTENNAMAXCUTCAR 25.643162 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.065 0.4 0.165 1.05 ;
        RECT 0.95 0.7 1.05 1.05 ;
        RECT 0.065 0.95 1.05 1.05 ;
      LAYER CUT01 ;
        RECT 0.07 0.45 0.16 0.54 ;
        RECT 0.955 0.74 1.045 0.83 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.117 LAYER MET1 ;
    ANTENNAMAXCUTCAR 51.286325 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.295 0.4 0.395 0.85 ;
        RECT 0.74 0.5 0.84 0.85 ;
        RECT 0.295 0.75 0.84 0.85 ;
        RECT 0.74 0.5 1.25 0.6 ;
        RECT 1.15 0.5 1.25 0.79 ;
        RECT 1.15 0.69 1.49 0.79 ;
        RECT 1.39 0.69 1.49 0.875 ;
      LAYER CUT01 ;
        RECT 0.3 0.45 0.39 0.54 ;
        RECT 0.645 0.755 0.735 0.845 ;
        RECT 1.395 0.735 1.485 0.825 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.51 1.24 0.61 1.96 ;
        RECT 1.03 1.4 1.13 1.96 ;
        RECT 1.575 1.26 1.675 1.96 ;
        RECT 2.11 1.26 2.21 1.96 ;
        RECT 2.63 1.24 2.73 1.96 ;
        RECT 0 1.64 2.8 1.96 ;
      LAYER CUT01 ;
        RECT 0.515 1.5 0.605 1.59 ;
        RECT 0.515 1.28 0.605 1.37 ;
        RECT 1.035 1.45 1.125 1.54 ;
        RECT 1.58 1.5 1.67 1.59 ;
        RECT 1.58 1.3 1.67 1.39 ;
        RECT 2.115 1.5 2.205 1.59 ;
        RECT 2.115 1.3 2.205 1.39 ;
        RECT 2.635 1.5 2.725 1.59 ;
        RECT 2.635 1.28 2.725 1.37 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.53 -0.16 0.63 0.55 ;
        RECT 1.55 -0.16 1.65 0.36 ;
        RECT 2.07 -0.16 2.25 0.32 ;
        RECT 2.63 -0.16 2.73 0.555 ;
        RECT 0 -0.16 2.8 0.16 ;
      LAYER CUT01 ;
        RECT 0.535 0.42 0.625 0.51 ;
        RECT 0.535 0.21 0.625 0.3 ;
        RECT 1.555 0.225 1.645 0.315 ;
        RECT 2.115 0.225 2.205 0.315 ;
        RECT 2.635 0.425 2.725 0.515 ;
        RECT 2.635 0.225 2.725 0.315 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4372 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 1.815 0.96 1.985 1.295 ;
        RECT 1.815 0.44 2.505 0.6 ;
        RECT 2.305 0.44 2.505 1.12 ;
        RECT 1.815 0.96 2.505 1.12 ;
        RECT 2.335 0.44 2.505 1.295 ;
      LAYER CUT01 ;
        RECT 1.855 1.195 1.945 1.285 ;
        RECT 1.855 0.975 1.945 1.065 ;
        RECT 1.855 0.47 1.945 0.56 ;
        RECT 2.375 1.195 2.465 1.285 ;
        RECT 2.375 0.975 2.465 1.065 ;
        RECT 2.375 0.47 2.465 0.56 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT -0.5 -0.5 3.3 0.78 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 3.3 2.3 ;
    END
  END VNW
  OBS
    LAYER MET1 ;
      RECT 0.99 0.31 1.45 0.41 ;
      RECT 1.35 0.31 1.45 0.575 ;
      RECT 1.35 0.475 1.69 0.575 ;
      RECT 1.59 0.72 2.165 0.82 ;
      RECT 1.59 0.475 1.69 1.1 ;
      RECT 1.29 1 1.69 1.1 ;
      RECT 0.73 1.15 1.39 1.25 ;
      RECT 1.29 1 1.39 1.385 ;
      RECT 0.77 1.15 0.87 1.485 ;
  END
END SC22ISOANDCLXL1

MACRO SC22ISOANDCLXP1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22ISOANDCLXP1 0 0 ;
  SIZE 4.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE CORE1800 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.1755 LAYER MET1 ;
    ANTENNAMAXCUTCAR 51.286325 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.065 0.4 0.165 1.05 ;
        RECT 0.955 0.7 1.055 1.05 ;
        RECT 1.915 0.69 2.015 1.05 ;
        RECT 0.065 0.95 2.015 1.05 ;
      LAYER CUT01 ;
        RECT 0.07 0.45 0.16 0.54 ;
        RECT 0.96 0.74 1.05 0.83 ;
        RECT 1.92 0.735 2.01 0.825 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.1755 LAYER MET1 ;
    ANTENNAMAXCUTCAR 51.286325 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.295 0.4 0.395 0.85 ;
        RECT 0.745 0.5 0.845 0.85 ;
        RECT 0.295 0.75 0.845 0.85 ;
        RECT 0.745 0.5 1.255 0.6 ;
        RECT 1.155 0.5 1.255 0.85 ;
        RECT 1.155 0.74 1.7 0.85 ;
      LAYER CUT01 ;
        RECT 0.3 0.45 0.39 0.54 ;
        RECT 0.65 0.755 0.74 0.845 ;
        RECT 1.56 0.74 1.65 0.83 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.515 1.24 0.615 1.96 ;
        RECT 1.035 1.4 1.135 1.96 ;
        RECT 1.555 1.4 1.655 1.96 ;
        RECT 2.1 1.4 2.2 1.96 ;
        RECT 2.645 1.25 2.745 1.96 ;
        RECT 3.165 1.24 3.265 1.96 ;
        RECT 3.685 1.24 3.785 1.96 ;
        RECT 4.205 1.24 4.305 1.96 ;
        RECT 0 1.64 4.4 1.96 ;
      LAYER CUT01 ;
        RECT 0.52 1.5 0.61 1.59 ;
        RECT 0.52 1.28 0.61 1.37 ;
        RECT 1.04 1.45 1.13 1.54 ;
        RECT 1.56 1.45 1.65 1.54 ;
        RECT 2.105 1.45 2.195 1.54 ;
        RECT 2.65 1.5 2.74 1.59 ;
        RECT 2.65 1.29 2.74 1.38 ;
        RECT 3.17 1.5 3.26 1.59 ;
        RECT 3.17 1.28 3.26 1.37 ;
        RECT 3.69 1.5 3.78 1.59 ;
        RECT 3.69 1.28 3.78 1.37 ;
        RECT 4.21 1.5 4.3 1.59 ;
        RECT 4.21 1.28 4.3 1.37 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.535 -0.16 0.635 0.55 ;
        RECT 1.555 -0.16 1.655 0.36 ;
        RECT 2.645 -0.16 2.745 0.57 ;
        RECT 3.165 -0.16 3.265 0.57 ;
        RECT 3.685 -0.16 3.785 0.57 ;
        RECT 4.205 -0.16 4.305 0.57 ;
        RECT 0 -0.16 4.4 0.16 ;
      LAYER CUT01 ;
        RECT 0.54 0.42 0.63 0.51 ;
        RECT 0.54 0.21 0.63 0.3 ;
        RECT 1.56 0.225 1.65 0.315 ;
        RECT 2.65 0.44 2.74 0.53 ;
        RECT 2.65 0.23 2.74 0.32 ;
        RECT 3.17 0.44 3.26 0.53 ;
        RECT 3.17 0.23 3.26 0.32 ;
        RECT 3.69 0.44 3.78 0.53 ;
        RECT 3.69 0.23 3.78 0.32 ;
        RECT 4.21 0.44 4.3 0.53 ;
        RECT 4.21 0.23 4.3 0.32 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.824 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 2.35 0.955 2.52 1.295 ;
        RECT 2.35 0.955 3.04 1.115 ;
        RECT 2.87 0.3 3.04 1.295 ;
        RECT 3.39 0.3 3.56 1.295 ;
        RECT 2.87 0.75 4.08 1.05 ;
        RECT 3.91 0.3 4.08 1.295 ;
      LAYER CUT01 ;
        RECT 2.39 1.195 2.48 1.285 ;
        RECT 2.39 0.975 2.48 1.065 ;
        RECT 2.91 1.195 3 1.285 ;
        RECT 2.91 0.975 3 1.065 ;
        RECT 2.91 0.505 3 0.595 ;
        RECT 2.91 0.305 3 0.395 ;
        RECT 3.43 1.195 3.52 1.285 ;
        RECT 3.43 0.975 3.52 1.065 ;
        RECT 3.43 0.505 3.52 0.595 ;
        RECT 3.43 0.305 3.52 0.395 ;
        RECT 3.95 1.195 4.04 1.285 ;
        RECT 3.95 0.975 4.04 1.065 ;
        RECT 3.95 0.505 4.04 0.595 ;
        RECT 3.95 0.305 4.04 0.395 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT -0.5 -0.5 4.9 0.78 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 4.9 2.3 ;
    END
  END VNW
  OBS
    LAYER MET1 ;
      RECT 0.995 0.31 1.455 0.41 ;
      RECT 1.355 0.31 1.455 0.575 ;
      RECT 1.355 0.475 2.22 0.575 ;
      RECT 2.12 0.715 2.73 0.815 ;
      RECT 2.12 0.475 2.22 1.25 ;
      RECT 0.735 1.15 2.22 1.25 ;
      RECT 0.775 1.15 0.875 1.485 ;
      RECT 1.295 1.15 1.395 1.485 ;
      RECT 1.815 1.15 1.915 1.485 ;
  END
END SC22ISOANDCLXP1

MACRO SC22ISOORCLXL1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22ISOORCLXL1 0 0 ;
  SIZE 3.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE CORE1800 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.13375 LAYER MET1 ;
    ANTENNAMAXCUTCAR 47.434535 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.82 0.4 0.92 0.85 ;
        RECT 0.82 0.55 1.7 0.65 ;
        RECT 1.6 0.55 1.7 0.8 ;
        RECT 1.6 0.7 1.975 0.8 ;
      LAYER CUT01 ;
        RECT 0.825 0.72 0.915 0.81 ;
        RECT 0.825 0.455 0.915 0.545 ;
        RECT 1.835 0.705 1.925 0.795 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.05725 LAYER MET1 ;
    ANTENNAMAXCUTCAR 52.406044 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.1 0.325 0.2 0.85 ;
        RECT 0.1 0.75 0.305 0.85 ;
        RECT 0.1 0.325 0.72 0.415 ;
      LAYER CUT01 ;
        RECT 0.165 0.755 0.255 0.845 ;
        RECT 0.58 0.325 0.67 0.415 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.345 1.25 0.445 1.96 ;
        RECT 1.315 1.4 1.415 1.96 ;
        RECT 2.17 1.25 2.27 1.96 ;
        RECT 2.69 1.26 2.79 1.96 ;
        RECT 3.21 1.24 3.31 1.96 ;
        RECT 0 1.64 3.4 1.96 ;
      LAYER CUT01 ;
        RECT 0.35 1.5 0.44 1.59 ;
        RECT 0.35 1.29 0.44 1.38 ;
        RECT 1.32 1.45 1.41 1.54 ;
        RECT 2.175 1.5 2.265 1.59 ;
        RECT 2.175 1.29 2.265 1.38 ;
        RECT 2.695 1.5 2.785 1.59 ;
        RECT 2.695 1.3 2.785 1.39 ;
        RECT 3.215 1.5 3.305 1.59 ;
        RECT 3.215 1.28 3.305 1.37 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.075 -0.16 0.175 0.225 ;
        RECT 1.055 -0.16 1.155 0.38 ;
        RECT 1.54 -0.16 1.72 0.23 ;
        RECT 2.105 -0.16 2.205 0.38 ;
        RECT 2.65 -0.16 2.83 0.32 ;
        RECT 3.21 -0.16 3.31 0.555 ;
        RECT 0 -0.16 3.4 0.16 ;
      LAYER CUT01 ;
        RECT 0.08 0.095 0.17 0.185 ;
        RECT 1.06 0.245 1.15 0.335 ;
        RECT 1.585 0.14 1.675 0.23 ;
        RECT 2.11 0.245 2.2 0.335 ;
        RECT 2.695 0.225 2.785 0.315 ;
        RECT 3.215 0.425 3.305 0.515 ;
        RECT 3.215 0.225 3.305 0.315 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4372 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 2.395 0.96 2.565 1.295 ;
        RECT 2.395 0.44 3.085 0.6 ;
        RECT 2.885 0.44 3.085 1.12 ;
        RECT 2.395 0.96 3.085 1.12 ;
        RECT 2.915 0.44 3.085 1.295 ;
      LAYER CUT01 ;
        RECT 2.435 1.195 2.525 1.285 ;
        RECT 2.435 0.975 2.525 1.065 ;
        RECT 2.435 0.47 2.525 0.56 ;
        RECT 2.955 1.195 3.045 1.285 ;
        RECT 2.955 0.975 3.045 1.065 ;
        RECT 2.955 0.47 3.045 0.56 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT -0.5 -0.5 3.9 0.78 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 3.9 2.3 ;
    END
  END VNW
  OBS
    LAYER MET1 ;
      RECT 0.3 0.505 0.55 0.605 ;
      RECT 1.27 0.75 1.46 0.85 ;
      RECT 0.45 0.505 0.55 1.05 ;
      RECT 1.27 0.75 1.37 1.05 ;
      RECT 0.08 0.95 1.37 1.05 ;
      RECT 0.08 0.95 0.18 1.325 ;
      RECT 1.275 0.35 1.985 0.45 ;
      RECT 1.885 0.35 1.985 0.59 ;
      RECT 1.885 0.49 2.2 0.59 ;
      RECT 2.1 0.72 2.745 0.82 ;
      RECT 2.1 0.49 2.2 1.05 ;
      RECT 1.845 0.95 2.2 1.05 ;
      RECT 0.795 1.15 1.945 1.25 ;
      RECT 1.845 0.95 1.945 1.39 ;
      RECT 0.835 1.15 0.935 1.485 ;
  END
END SC22ISOORCLXL1

MACRO SC22ISOORCLXP1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22ISOORCLXP1 0 0 ;
  SIZE 5.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE CORE1800 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.22275 LAYER MET1 ;
    ANTENNAMAXCUTCAR 59.118062 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.795 0.455 0.895 0.85 ;
        RECT 1.81 0.55 1.91 0.83 ;
        RECT 0.795 0.55 2.52 0.65 ;
        RECT 2.42 0.55 2.52 0.785 ;
        RECT 2.42 0.685 2.72 0.785 ;
        RECT 2.62 0.685 2.72 0.875 ;
      LAYER CUT01 ;
        RECT 0.8 0.72 0.89 0.81 ;
        RECT 0.8 0.5 0.89 0.59 ;
        RECT 1.815 0.69 1.905 0.78 ;
        RECT 2.625 0.735 2.715 0.825 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.05725 LAYER MET1 ;
    ANTENNAMAXCUTCAR 52.406044 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.09 0.32 0.19 0.85 ;
        RECT 0.09 0.75 0.3 0.85 ;
        RECT 0.09 0.32 0.71 0.41 ;
      LAYER CUT01 ;
        RECT 0.155 0.755 0.245 0.845 ;
        RECT 0.57 0.32 0.66 0.41 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.335 1.25 0.435 1.96 ;
        RECT 1.29 1.4 1.39 1.96 ;
        RECT 2.26 1.4 2.36 1.96 ;
        RECT 2.95 1.25 3.05 1.96 ;
        RECT 3.47 1.25 3.57 1.96 ;
        RECT 3.99 1.24 4.09 1.96 ;
        RECT 4.51 1.24 4.61 1.96 ;
        RECT 5.03 1.24 5.13 1.96 ;
        RECT 0 1.64 5.2 1.96 ;
      LAYER CUT01 ;
        RECT 0.34 1.5 0.43 1.59 ;
        RECT 0.34 1.29 0.43 1.38 ;
        RECT 1.295 1.45 1.385 1.54 ;
        RECT 2.265 1.45 2.355 1.54 ;
        RECT 2.955 1.5 3.045 1.59 ;
        RECT 2.955 1.29 3.045 1.38 ;
        RECT 3.475 1.5 3.565 1.59 ;
        RECT 3.475 1.29 3.565 1.38 ;
        RECT 3.995 1.5 4.085 1.59 ;
        RECT 3.995 1.28 4.085 1.37 ;
        RECT 4.515 1.5 4.605 1.59 ;
        RECT 4.515 1.28 4.605 1.37 ;
        RECT 5.035 1.5 5.125 1.59 ;
        RECT 5.035 1.28 5.125 1.37 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.065 -0.16 0.165 0.225 ;
        RECT 1.03 -0.16 1.13 0.375 ;
        RECT 1.515 -0.16 1.695 0.23 ;
        RECT 2.13 -0.16 2.31 0.23 ;
        RECT 2.82 -0.16 2.92 0.375 ;
        RECT 3.47 -0.16 3.57 0.57 ;
        RECT 3.99 -0.16 4.09 0.57 ;
        RECT 4.51 -0.16 4.61 0.57 ;
        RECT 5.03 -0.16 5.13 0.57 ;
        RECT 0 -0.16 5.2 0.16 ;
      LAYER CUT01 ;
        RECT 0.07 0.095 0.16 0.185 ;
        RECT 1.035 0.24 1.125 0.33 ;
        RECT 1.56 0.14 1.65 0.23 ;
        RECT 2.175 0.14 2.265 0.23 ;
        RECT 2.825 0.24 2.915 0.33 ;
        RECT 3.475 0.44 3.565 0.53 ;
        RECT 3.475 0.23 3.565 0.32 ;
        RECT 3.995 0.44 4.085 0.53 ;
        RECT 3.995 0.23 4.085 0.32 ;
        RECT 4.515 0.44 4.605 0.53 ;
        RECT 4.515 0.23 4.605 0.32 ;
        RECT 5.035 0.44 5.125 0.53 ;
        RECT 5.035 0.23 5.125 0.32 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.824 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 3.175 0.955 3.345 1.295 ;
        RECT 3.175 0.955 3.865 1.115 ;
        RECT 3.695 0.3 3.865 1.295 ;
        RECT 4.215 0.3 4.385 1.295 ;
        RECT 3.695 0.75 4.905 1.05 ;
        RECT 4.735 0.3 4.905 1.295 ;
      LAYER CUT01 ;
        RECT 3.215 1.195 3.305 1.285 ;
        RECT 3.215 0.975 3.305 1.065 ;
        RECT 3.735 1.195 3.825 1.285 ;
        RECT 3.735 0.975 3.825 1.065 ;
        RECT 3.735 0.505 3.825 0.595 ;
        RECT 3.735 0.305 3.825 0.395 ;
        RECT 4.255 1.195 4.345 1.285 ;
        RECT 4.255 0.975 4.345 1.065 ;
        RECT 4.255 0.505 4.345 0.595 ;
        RECT 4.255 0.305 4.345 0.395 ;
        RECT 4.775 1.195 4.865 1.285 ;
        RECT 4.775 0.975 4.865 1.065 ;
        RECT 4.775 0.505 4.865 0.595 ;
        RECT 4.775 0.305 4.865 0.395 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT -0.5 -0.5 5.7 0.78 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 5.7 2.3 ;
    END
  END VNW
  OBS
    LAYER MET1 ;
      RECT 0.29 0.505 0.54 0.605 ;
      RECT 1.245 0.75 1.435 0.85 ;
      RECT 2.1 0.75 2.32 0.85 ;
      RECT 0.44 0.505 0.54 1.05 ;
      RECT 1.29 0.75 1.39 1.05 ;
      RECT 2.1 0.75 2.2 1.05 ;
      RECT 0.07 0.95 2.2 1.05 ;
      RECT 0.07 0.95 0.17 1.325 ;
      RECT 1.25 0.35 2.72 0.45 ;
      RECT 2.62 0.35 2.72 0.585 ;
      RECT 2.62 0.485 2.94 0.585 ;
      RECT 2.84 0.715 3.555 0.815 ;
      RECT 2.84 0.485 2.94 1.11 ;
      RECT 2.72 1.01 2.94 1.11 ;
      RECT 0.775 1.15 2.82 1.25 ;
      RECT 2.72 1.01 2.82 1.44 ;
      RECT 0.815 1.15 0.915 1.485 ;
      RECT 1.8 1.15 1.9 1.485 ;
  END
END SC22ISOORCLXP1

MACRO SC22LSBIANDCLXL1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSBIANDCLXL1 0 0 ;
  SIZE 5.6 BY 3.6 ;
  SYMMETRY X Y ;
  SITE WCORE3600 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.0585 LAYER MET1 ;
    ANTENNAMAXCUTCAR 51.286325 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VYY ;
    PORT
      LAYER MET1 ;
        RECT 1.3 0.4 1.4 0.85 ;
        RECT 1.3 0.74 1.81 0.85 ;
      LAYER CUT01 ;
        RECT 1.305 0.45 1.395 0.54 ;
        RECT 1.675 0.745 1.765 0.835 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.0585 LAYER MET1 ;
    ANTENNAMAXCUTCAR 51.286325 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 5.15 0.4 5.25 1.225 ;
        RECT 5.15 1.125 5.47 1.225 ;
      LAYER CUT01 ;
        RECT 5.155 0.45 5.245 0.54 ;
        RECT 5.335 1.13 5.425 1.22 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 0.5 2.82 ;
        RECT 3.5 0.78 6.1 2.82 ;
      LAYER MET1 ;
        RECT 3.61 1.595 3.79 1.96 ;
        RECT 4.13 1.64 4.31 2.005 ;
        RECT 4.19 1.595 4.37 1.96 ;
        RECT 4.78 1.595 4.96 1.96 ;
        RECT 5.09 1.595 5.27 1.96 ;
        RECT 5.12 1.64 5.3 2.005 ;
        RECT 0 1.64 5.6 1.96 ;
      LAYER CUT01 ;
        RECT 0.175 1.86 0.265 1.95 ;
        RECT 0.175 1.65 0.265 1.74 ;
        RECT 3.655 1.595 3.745 1.685 ;
        RECT 4.175 1.915 4.265 2.005 ;
        RECT 4.235 1.595 4.325 1.685 ;
        RECT 4.825 1.595 4.915 1.685 ;
        RECT 5.135 1.595 5.225 1.685 ;
        RECT 5.165 1.915 5.255 2.005 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 1.965 3.065 2.065 3.76 ;
        RECT 5.43 3.245 5.53 3.76 ;
        RECT 0 3.44 5.6 3.76 ;
        RECT 1.65 -0.16 1.75 0.535 ;
        RECT 3.675 -0.16 3.775 0.56 ;
        RECT 4.23 -0.16 4.33 0.56 ;
        RECT 0 -0.16 5.6 0.16 ;
      LAYER CUT01 ;
        RECT 1.655 0.405 1.745 0.495 ;
        RECT 1.655 0.205 1.745 0.295 ;
        RECT 1.97 3.305 2.06 3.395 ;
        RECT 1.97 3.105 2.06 3.195 ;
        RECT 3.68 0.43 3.77 0.52 ;
        RECT 3.68 0.23 3.77 0.32 ;
        RECT 4.235 0.43 4.325 0.52 ;
        RECT 4.235 0.23 4.325 0.32 ;
        RECT 5.435 3.295 5.525 3.385 ;
    END
  END VSS
  PIN VYY
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT 1.5 0.78 2.5 2.82 ;
      LAYER MET1 ;
        RECT 1.65 2.125 1.75 2.46 ;
        RECT 1.965 2.125 2.065 2.46 ;
        RECT 0.06 2.125 5.54 2.275 ;
        RECT 1.65 1.14 1.75 1.475 ;
        RECT 0.06 1.325 5.54 1.475 ;
      LAYER CUT01 ;
        RECT 1.655 2.33 1.745 2.42 ;
        RECT 1.655 2.13 1.745 2.22 ;
        RECT 1.655 1.38 1.745 1.47 ;
        RECT 1.655 1.18 1.745 1.27 ;
        RECT 1.97 2.33 2.06 2.42 ;
        RECT 1.97 2.13 2.06 2.22 ;
    END
  END VYY
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4477 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 3.9 0.3 4.07 1.185 ;
        RECT 3.9 0.7 4.66 0.9 ;
        RECT 4.49 0.3 4.66 1.185 ;
      LAYER CUT01 ;
        RECT 3.94 1.075 4.03 1.165 ;
        RECT 3.94 0.505 4.03 0.595 ;
        RECT 3.94 0.305 4.03 0.395 ;
        RECT 4.53 1.075 4.62 1.165 ;
        RECT 4.53 0.505 4.62 0.595 ;
        RECT 4.53 0.305 4.62 0.395 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT 0.5 -0.5 1.5 4.1 ;
        RECT 2.5 -0.5 3.5 4.1 ;
        RECT -0.5 -0.5 6.1 0.78 ;
        RECT -0.5 2.82 6.1 4.1 ;
    END
  END VPW
  OBS
    LAYER MET1 ;
      RECT 1.91 0.385 2.36 0.485 ;
      RECT 1.91 0.285 2.01 1.225 ;
      RECT 1.865 1.125 3.575 1.225 ;
      RECT 2.18 2.375 2.37 2.475 ;
      RECT 4.54 2.77 4.805 2.87 ;
      RECT 4.54 2.77 4.64 3.075 ;
      RECT 4.055 2.975 4.64 3.075 ;
      RECT 4.055 2.975 4.155 3.28 ;
      RECT 2.225 3.18 4.155 3.28 ;
      RECT 2.225 2.375 2.325 3.315 ;
      RECT 3.52 2.375 3.815 2.475 ;
      RECT 4.33 2.575 5.145 2.675 ;
      RECT 4.33 2.575 4.43 2.875 ;
      RECT 3.855 2.775 4.43 2.875 ;
      RECT 5.045 2.575 5.145 2.89 ;
      RECT 3.52 2.375 3.62 3.085 ;
      RECT 3.855 2.775 3.955 3.085 ;
      RECT 3.52 2.985 3.955 3.085 ;
      RECT 4.255 3.19 5.31 3.29 ;
      RECT 4.005 2.375 5.53 2.475 ;
      RECT 4.005 2.375 4.105 2.675 ;
      RECT 3.72 2.575 4.105 2.675 ;
      RECT 5.43 2.375 5.53 3.09 ;
      RECT 4.755 2.99 5.53 3.09 ;
  END
END SC22LSBIANDCLXL1

MACRO SC22LSBIANDCLXP1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSBIANDCLXP1 0 0 ;
  SIZE 7.2 BY 3.6 ;
  SYMMETRY X Y ;
  SITE WCORE3600 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.117 LAYER MET1 ;
    ANTENNAMAXCUTCAR 25.643162 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VYY ;
    PORT
      LAYER MET1 ;
        RECT 1.3 0.4 1.4 0.85 ;
        RECT 1.3 0.74 1.81 0.85 ;
      LAYER CUT01 ;
        RECT 1.305 0.45 1.395 0.54 ;
        RECT 1.675 0.745 1.765 0.835 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.117 LAYER MET1 ;
    ANTENNAMAXCUTCAR 32.00256 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 6.55 0.4 6.65 1.225 ;
        RECT 6.505 1.125 6.695 1.225 ;
      LAYER CUT01 ;
        RECT 6.555 1.13 6.645 1.22 ;
        RECT 6.555 0.45 6.645 0.54 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 0.5 2.82 ;
        RECT 3.7 0.78 7.7 2.82 ;
      LAYER MET1 ;
        RECT 3.81 1.595 3.99 1.96 ;
        RECT 4.33 1.64 4.51 2.005 ;
        RECT 4.4 1.595 4.58 1.96 ;
        RECT 4.99 1.595 5.17 1.96 ;
        RECT 5.32 1.64 5.5 2.005 ;
        RECT 5.58 1.595 5.76 1.96 ;
        RECT 6.17 1.595 6.35 1.96 ;
        RECT 6.31 1.64 6.49 2.005 ;
        RECT 6.9 1.64 7.08 2.005 ;
        RECT 6.915 1.595 7.095 1.96 ;
        RECT 0 1.64 7.2 1.96 ;
      LAYER CUT01 ;
        RECT 0.175 1.86 0.265 1.95 ;
        RECT 0.175 1.65 0.265 1.74 ;
        RECT 3.855 1.595 3.945 1.685 ;
        RECT 4.375 1.915 4.465 2.005 ;
        RECT 4.445 1.595 4.535 1.685 ;
        RECT 5.035 1.595 5.125 1.685 ;
        RECT 5.365 1.915 5.455 2.005 ;
        RECT 5.625 1.595 5.715 1.685 ;
        RECT 6.215 1.595 6.305 1.685 ;
        RECT 6.355 1.915 6.445 2.005 ;
        RECT 6.945 1.915 7.035 2.005 ;
        RECT 6.96 1.595 7.05 1.685 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 1.93 3.065 2.03 3.76 ;
        RECT 2.45 3.065 2.55 3.76 ;
        RECT 6.31 3.41 6.49 3.76 ;
        RECT 6.905 3.065 7.005 3.76 ;
        RECT 0 3.44 7.2 3.76 ;
        RECT 1.65 -0.16 1.75 0.535 ;
        RECT 2.17 -0.16 2.27 0.535 ;
        RECT 3.885 -0.16 3.985 0.56 ;
        RECT 4.44 -0.16 4.54 0.56 ;
        RECT 5.03 -0.16 5.13 0.56 ;
        RECT 5.585 -0.16 5.685 0.56 ;
        RECT 0 -0.16 7.2 0.16 ;
      LAYER CUT01 ;
        RECT 1.655 0.405 1.745 0.495 ;
        RECT 1.655 0.205 1.745 0.295 ;
        RECT 1.935 3.305 2.025 3.395 ;
        RECT 1.935 3.105 2.025 3.195 ;
        RECT 2.175 0.405 2.265 0.495 ;
        RECT 2.175 0.205 2.265 0.295 ;
        RECT 2.455 3.305 2.545 3.395 ;
        RECT 2.455 3.105 2.545 3.195 ;
        RECT 3.89 0.43 3.98 0.52 ;
        RECT 3.89 0.23 3.98 0.32 ;
        RECT 4.445 0.43 4.535 0.52 ;
        RECT 4.445 0.23 4.535 0.32 ;
        RECT 5.035 0.43 5.125 0.52 ;
        RECT 5.035 0.23 5.125 0.32 ;
        RECT 5.59 0.43 5.68 0.52 ;
        RECT 5.59 0.23 5.68 0.32 ;
        RECT 6.355 3.41 6.445 3.5 ;
        RECT 6.91 3.305 7 3.395 ;
        RECT 6.91 3.105 7 3.195 ;
    END
  END VSS
  PIN VYY
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT 1.5 0.78 2.7 2.82 ;
      LAYER MET1 ;
        RECT 1.65 2.125 1.75 2.46 ;
        RECT 1.93 2.125 2.03 2.46 ;
        RECT 2.45 2.125 2.55 2.46 ;
        RECT 0.06 2.125 7.14 2.275 ;
        RECT 1.65 1.14 1.75 1.475 ;
        RECT 2.17 1.14 2.27 1.475 ;
        RECT 0.06 1.325 7.14 1.475 ;
      LAYER CUT01 ;
        RECT 1.655 2.33 1.745 2.42 ;
        RECT 1.655 2.13 1.745 2.22 ;
        RECT 1.655 1.38 1.745 1.47 ;
        RECT 1.655 1.18 1.745 1.27 ;
        RECT 1.935 2.33 2.025 2.42 ;
        RECT 1.935 2.13 2.025 2.22 ;
        RECT 2.175 1.38 2.265 1.47 ;
        RECT 2.175 1.18 2.265 1.27 ;
        RECT 2.455 2.33 2.545 2.42 ;
        RECT 2.455 2.13 2.545 2.22 ;
    END
  END VYY
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.824 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 4.11 0.3 4.28 1.185 ;
        RECT 4.7 0.3 4.87 1.185 ;
        RECT 5.29 0.3 5.46 1.185 ;
        RECT 4.11 0.75 6.05 1.05 ;
        RECT 5.88 0.75 6.05 1.185 ;
      LAYER CUT01 ;
        RECT 4.15 1.075 4.24 1.165 ;
        RECT 4.15 0.505 4.24 0.595 ;
        RECT 4.15 0.305 4.24 0.395 ;
        RECT 4.74 1.075 4.83 1.165 ;
        RECT 4.74 0.505 4.83 0.595 ;
        RECT 4.74 0.305 4.83 0.395 ;
        RECT 5.33 1.075 5.42 1.165 ;
        RECT 5.33 0.505 5.42 0.595 ;
        RECT 5.33 0.305 5.42 0.395 ;
        RECT 5.92 1.075 6.01 1.165 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT 0.5 -0.5 1.5 4.1 ;
        RECT 2.7 -0.5 3.7 4.1 ;
        RECT -0.5 -0.5 7.7 0.78 ;
        RECT -0.5 2.82 7.7 4.1 ;
    END
  END VPW
  OBS
    LAYER MET1 ;
      RECT 1.91 0.785 2.63 0.885 ;
      RECT 1.91 0.285 2.01 1.225 ;
      RECT 2.53 0.4 2.63 1.225 ;
      RECT 1.865 1.125 2.055 1.225 ;
      RECT 2.53 1.125 2.815 1.225 ;
      RECT 2.145 2.375 2.335 2.475 ;
      RECT 4.825 2.775 5.005 2.875 ;
      RECT 5.605 2.775 6 2.875 ;
      RECT 2.19 2.8 2.87 2.9 ;
      RECT 4.865 2.775 4.965 3.075 ;
      RECT 5.605 2.775 5.705 3.075 ;
      RECT 4.32 2.975 5.705 3.075 ;
      RECT 2.77 2.8 2.87 3.28 ;
      RECT 4.32 2.975 4.42 3.28 ;
      RECT 2.77 3.18 4.42 3.28 ;
      RECT 2.19 2.375 2.29 3.315 ;
      RECT 3.44 2.375 4.015 2.475 ;
      RECT 4.54 2.575 6.335 2.675 ;
      RECT 5.355 2.575 5.455 2.875 ;
      RECT 4.54 2.575 4.64 2.875 ;
      RECT 4.12 2.775 4.64 2.875 ;
      RECT 5.315 2.775 5.495 2.875 ;
      RECT 6.235 2.575 6.335 2.89 ;
      RECT 3.44 2.375 3.54 3.08 ;
      RECT 4.12 2.775 4.22 3.08 ;
      RECT 3.44 2.98 4.22 3.08 ;
      RECT 4.205 2.375 6.745 2.475 ;
      RECT 4.205 2.375 4.305 2.675 ;
      RECT 3.64 2.575 4.305 2.675 ;
      RECT 6.645 2.375 6.745 3.09 ;
      RECT 5.815 2.99 6.745 3.09 ;
      RECT 4.52 3.19 6.785 3.29 ;
  END
END SC22LSBIANDCLXP1

MACRO SC22LSBICLXL1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSBICLXL1 0 0 ;
  SIZE 5.4 BY 3.6 ;
  SYMMETRY X Y ;
  SITE WCORE3600 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.0585 LAYER MET1 ;
    ANTENNAMAXCUTCAR 51.286325 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VYY ;
    PORT
      LAYER MET1 ;
        RECT 1.3 0.4 1.4 0.85 ;
        RECT 1.3 0.74 1.81 0.85 ;
      LAYER CUT01 ;
        RECT 1.305 0.45 1.395 0.54 ;
        RECT 1.675 0.745 1.765 0.835 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 0.5 2.82 ;
        RECT 3.5 0.78 5.9 2.82 ;
      LAYER MET1 ;
        RECT 3.61 1.595 3.79 1.96 ;
        RECT 4.14 1.64 4.32 2.005 ;
        RECT 4.2 1.595 4.38 1.96 ;
        RECT 4.79 1.595 4.97 1.96 ;
        RECT 5.115 1.595 5.295 1.96 ;
        RECT 5.13 1.64 5.31 2.005 ;
        RECT 0 1.64 5.4 1.96 ;
      LAYER CUT01 ;
        RECT 0.175 1.86 0.265 1.95 ;
        RECT 0.175 1.65 0.265 1.74 ;
        RECT 3.655 1.595 3.745 1.685 ;
        RECT 4.185 1.915 4.275 2.005 ;
        RECT 4.245 1.595 4.335 1.685 ;
        RECT 4.835 1.595 4.925 1.685 ;
        RECT 5.16 1.595 5.25 1.685 ;
        RECT 5.175 1.915 5.265 2.005 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 1.965 3.065 2.065 3.76 ;
        RECT 4.35 3.2 4.45 3.76 ;
        RECT 0 3.44 5.4 3.76 ;
        RECT 1.65 -0.16 1.75 0.535 ;
        RECT 3.685 -0.16 3.785 0.56 ;
        RECT 4.24 -0.16 4.34 0.56 ;
        RECT 0 -0.16 5.4 0.16 ;
      LAYER CUT01 ;
        RECT 1.655 0.405 1.745 0.495 ;
        RECT 1.655 0.205 1.745 0.295 ;
        RECT 1.97 3.305 2.06 3.395 ;
        RECT 1.97 3.105 2.06 3.195 ;
        RECT 3.69 0.43 3.78 0.52 ;
        RECT 3.69 0.23 3.78 0.32 ;
        RECT 4.245 0.43 4.335 0.52 ;
        RECT 4.245 0.23 4.335 0.32 ;
        RECT 4.355 3.245 4.445 3.335 ;
    END
  END VSS
  PIN VYY
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT 1.5 0.78 2.5 2.82 ;
      LAYER MET1 ;
        RECT 1.65 2.125 1.75 2.46 ;
        RECT 1.965 2.125 2.065 2.46 ;
        RECT 0.06 2.125 5.34 2.275 ;
        RECT 1.65 1.14 1.75 1.475 ;
        RECT 0.06 1.325 5.34 1.475 ;
      LAYER CUT01 ;
        RECT 1.655 2.33 1.745 2.42 ;
        RECT 1.655 2.13 1.745 2.22 ;
        RECT 1.655 1.38 1.745 1.47 ;
        RECT 1.655 1.18 1.745 1.27 ;
        RECT 1.97 2.33 2.06 2.42 ;
        RECT 1.97 2.13 2.06 2.22 ;
    END
  END VYY
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4477 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 3.91 0.3 4.08 1.185 ;
        RECT 3.91 0.7 4.67 0.9 ;
        RECT 4.5 0.3 4.67 1.185 ;
      LAYER CUT01 ;
        RECT 3.95 1.075 4.04 1.165 ;
        RECT 3.95 0.505 4.04 0.595 ;
        RECT 3.95 0.305 4.04 0.395 ;
        RECT 4.54 1.075 4.63 1.165 ;
        RECT 4.54 0.505 4.63 0.595 ;
        RECT 4.54 0.305 4.63 0.395 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT 0.5 -0.5 1.5 4.1 ;
        RECT 2.5 -0.5 3.5 4.1 ;
        RECT -0.5 -0.5 5.9 0.78 ;
        RECT -0.5 2.82 5.9 4.1 ;
    END
  END VPW
  OBS
    LAYER MET1 ;
      RECT 1.91 0.385 2.36 0.485 ;
      RECT 1.91 0.285 2.01 1.225 ;
      RECT 1.865 1.125 3.575 1.225 ;
      RECT 2.18 2.375 2.37 2.475 ;
      RECT 4.57 2.77 4.8 2.87 ;
      RECT 4.57 2.77 4.67 3.075 ;
      RECT 4.14 2.975 4.67 3.075 ;
      RECT 4.14 2.975 4.24 3.28 ;
      RECT 2.225 3.18 4.24 3.28 ;
      RECT 2.225 2.375 2.325 3.315 ;
      RECT 3.53 2.375 3.825 2.475 ;
      RECT 4.35 2.575 5.135 2.675 ;
      RECT 4.35 2.575 4.45 2.875 ;
      RECT 3.93 2.775 4.45 2.875 ;
      RECT 5.035 2.575 5.135 2.925 ;
      RECT 3.53 2.375 3.63 3.08 ;
      RECT 3.93 2.775 4.03 3.08 ;
      RECT 3.53 2.98 4.03 3.08 ;
      RECT 4.015 2.375 5.335 2.475 ;
      RECT 4.015 2.375 4.115 2.675 ;
      RECT 3.73 2.575 4.115 2.675 ;
      RECT 5.235 2.375 5.335 3.275 ;
      RECT 4.635 3.175 5.335 3.275 ;
  END
END SC22LSBICLXL1

MACRO SC22LSBICLXP1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSBICLXP1 0 0 ;
  SIZE 6.6 BY 3.6 ;
  SYMMETRY X Y ;
  SITE WCORE3600 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.117 LAYER MET1 ;
    ANTENNAMAXCUTCAR 25.643162 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VYY ;
    PORT
      LAYER MET1 ;
        RECT 1.3 0.4 1.4 0.85 ;
        RECT 1.3 0.74 1.81 0.85 ;
      LAYER CUT01 ;
        RECT 1.305 0.45 1.395 0.54 ;
        RECT 1.675 0.745 1.765 0.835 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 0.5 2.82 ;
        RECT 3.7 0.78 7.1 2.82 ;
      LAYER MET1 ;
        RECT 3.81 1.595 3.99 1.96 ;
        RECT 3.935 1.64 4.115 2.005 ;
        RECT 4.34 1.64 4.52 2.005 ;
        RECT 4.4 1.595 4.58 1.96 ;
        RECT 4.99 1.595 5.17 1.96 ;
        RECT 5.33 1.64 5.51 2.005 ;
        RECT 5.58 1.595 5.76 1.96 ;
        RECT 6.17 1.595 6.35 1.96 ;
        RECT 6.32 1.64 6.5 2.005 ;
        RECT 0 1.64 6.6 1.96 ;
      LAYER CUT01 ;
        RECT 0.175 1.86 0.265 1.95 ;
        RECT 0.175 1.65 0.265 1.74 ;
        RECT 3.855 1.595 3.945 1.685 ;
        RECT 3.98 1.915 4.07 2.005 ;
        RECT 4.385 1.915 4.475 2.005 ;
        RECT 4.445 1.595 4.535 1.685 ;
        RECT 5.035 1.595 5.125 1.685 ;
        RECT 5.375 1.915 5.465 2.005 ;
        RECT 5.625 1.595 5.715 1.685 ;
        RECT 6.215 1.595 6.305 1.685 ;
        RECT 6.365 1.915 6.455 2.005 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 1.93 3.065 2.03 3.76 ;
        RECT 2.45 3.065 2.55 3.76 ;
        RECT 4.53 3.25 4.63 3.76 ;
        RECT 5.605 3.25 5.705 3.76 ;
        RECT 6.125 3.25 6.225 3.76 ;
        RECT 0 3.44 6.6 3.76 ;
        RECT 1.65 -0.16 1.75 0.535 ;
        RECT 2.17 -0.16 2.27 0.535 ;
        RECT 3.885 -0.16 3.985 0.56 ;
        RECT 4.44 -0.16 4.54 0.56 ;
        RECT 5.03 -0.16 5.13 0.56 ;
        RECT 5.585 -0.16 5.685 0.56 ;
        RECT 0 -0.16 6.6 0.16 ;
      LAYER CUT01 ;
        RECT 1.655 0.405 1.745 0.495 ;
        RECT 1.655 0.205 1.745 0.295 ;
        RECT 1.935 3.305 2.025 3.395 ;
        RECT 1.935 3.105 2.025 3.195 ;
        RECT 2.175 0.405 2.265 0.495 ;
        RECT 2.175 0.205 2.265 0.295 ;
        RECT 2.455 3.305 2.545 3.395 ;
        RECT 2.455 3.105 2.545 3.195 ;
        RECT 3.89 0.43 3.98 0.52 ;
        RECT 3.89 0.23 3.98 0.32 ;
        RECT 4.445 0.43 4.535 0.52 ;
        RECT 4.445 0.23 4.535 0.32 ;
        RECT 4.535 3.295 4.625 3.385 ;
        RECT 5.035 0.43 5.125 0.52 ;
        RECT 5.035 0.23 5.125 0.32 ;
        RECT 5.59 0.43 5.68 0.52 ;
        RECT 5.59 0.23 5.68 0.32 ;
        RECT 5.61 3.295 5.7 3.385 ;
        RECT 6.13 3.295 6.22 3.385 ;
    END
  END VSS
  PIN VYY
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT 1.5 0.78 2.7 2.82 ;
      LAYER MET1 ;
        RECT 1.65 2.125 1.75 2.46 ;
        RECT 1.93 2.125 2.03 2.46 ;
        RECT 2.45 2.125 2.55 2.46 ;
        RECT 0.06 2.125 6.54 2.275 ;
        RECT 1.65 1.14 1.75 1.475 ;
        RECT 2.17 1.14 2.27 1.475 ;
        RECT 0.06 1.325 6.54 1.475 ;
      LAYER CUT01 ;
        RECT 1.655 2.33 1.745 2.42 ;
        RECT 1.655 2.13 1.745 2.22 ;
        RECT 1.655 1.38 1.745 1.47 ;
        RECT 1.655 1.18 1.745 1.27 ;
        RECT 1.935 2.33 2.025 2.42 ;
        RECT 1.935 2.13 2.025 2.22 ;
        RECT 2.175 1.38 2.265 1.47 ;
        RECT 2.175 1.18 2.265 1.27 ;
        RECT 2.455 2.33 2.545 2.42 ;
        RECT 2.455 2.13 2.545 2.22 ;
    END
  END VYY
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.824 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 4.11 0.3 4.28 1.185 ;
        RECT 4.7 0.3 4.87 1.185 ;
        RECT 5.29 0.3 5.46 1.185 ;
        RECT 4.11 0.75 6.05 1.05 ;
        RECT 5.88 0.75 6.05 1.185 ;
      LAYER CUT01 ;
        RECT 4.15 1.075 4.24 1.165 ;
        RECT 4.15 0.505 4.24 0.595 ;
        RECT 4.15 0.305 4.24 0.395 ;
        RECT 4.74 1.075 4.83 1.165 ;
        RECT 4.74 0.505 4.83 0.595 ;
        RECT 4.74 0.305 4.83 0.395 ;
        RECT 5.33 1.075 5.42 1.165 ;
        RECT 5.33 0.505 5.42 0.595 ;
        RECT 5.33 0.305 5.42 0.395 ;
        RECT 5.92 1.075 6.01 1.165 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT 0.5 -0.5 1.5 4.1 ;
        RECT 2.7 -0.5 3.7 4.1 ;
        RECT -0.5 -0.5 7.1 0.78 ;
        RECT -0.5 2.82 7.1 4.1 ;
    END
  END VPW
  OBS
    LAYER MET1 ;
      RECT 1.91 0.785 2.63 0.885 ;
      RECT 1.91 0.285 2.01 1.225 ;
      RECT 2.53 0.4 2.63 1.225 ;
      RECT 1.865 1.125 2.055 1.225 ;
      RECT 2.53 1.125 2.815 1.225 ;
      RECT 2.145 2.375 2.335 2.475 ;
      RECT 4.835 2.775 5.015 2.875 ;
      RECT 5.615 2.775 6.01 2.875 ;
      RECT 2.19 2.8 2.87 2.9 ;
      RECT 4.875 2.775 4.975 3.075 ;
      RECT 5.615 2.775 5.715 3.075 ;
      RECT 4.33 2.975 5.715 3.075 ;
      RECT 2.77 2.8 2.87 3.28 ;
      RECT 4.33 2.975 4.43 3.28 ;
      RECT 2.77 3.18 4.43 3.28 ;
      RECT 2.19 2.375 2.29 3.315 ;
      RECT 3.44 2.375 4.025 2.475 ;
      RECT 4.55 2.575 6.325 2.675 ;
      RECT 5.365 2.575 5.465 2.875 ;
      RECT 4.55 2.575 4.65 2.875 ;
      RECT 4.13 2.775 4.65 2.875 ;
      RECT 5.325 2.775 5.505 2.875 ;
      RECT 6.225 2.575 6.325 2.91 ;
      RECT 3.44 2.375 3.54 3.08 ;
      RECT 4.13 2.775 4.23 3.08 ;
      RECT 3.44 2.98 4.23 3.08 ;
      RECT 4.215 2.375 6.525 2.475 ;
      RECT 4.215 2.375 4.315 2.675 ;
      RECT 3.64 2.575 4.315 2.675 ;
      RECT 6.425 2.375 6.525 3.13 ;
      RECT 5.825 3.03 6.525 3.13 ;
  END
END SC22LSBICLXP1

MACRO SC22LSBIORCLXL1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSBIORCLXL1 0 0 ;
  SIZE 5.8 BY 3.6 ;
  SYMMETRY X Y ;
  SITE WCORE3600 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.0585 LAYER MET1 ;
    ANTENNAMAXCUTCAR 51.286325 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VYY ;
    PORT
      LAYER MET1 ;
        RECT 1.3 0.4 1.4 0.85 ;
        RECT 1.3 0.74 1.81 0.85 ;
      LAYER CUT01 ;
        RECT 1.305 0.45 1.395 0.54 ;
        RECT 1.675 0.745 1.765 0.835 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.0585 LAYER MET1 ;
    ANTENNAMAXCUTCAR 51.286325 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 5.4 0.4 5.5 0.85 ;
        RECT 5.065 0.74 5.5 0.85 ;
      LAYER CUT01 ;
        RECT 5.11 0.745 5.2 0.835 ;
        RECT 5.405 0.45 5.495 0.54 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 0.5 2.82 ;
        RECT 3.5 0.78 6.3 2.82 ;
      LAYER MET1 ;
        RECT 3.61 1.595 3.79 1.96 ;
        RECT 4.2 1.595 4.38 1.96 ;
        RECT 4.79 1.595 4.97 1.96 ;
        RECT 5.325 1.64 5.505 2.005 ;
        RECT 5.51 1.595 5.69 1.96 ;
        RECT 0 1.64 5.8 1.96 ;
      LAYER CUT01 ;
        RECT 0.175 1.86 0.265 1.95 ;
        RECT 0.175 1.65 0.265 1.74 ;
        RECT 3.655 1.595 3.745 1.685 ;
        RECT 4.245 1.595 4.335 1.685 ;
        RECT 4.835 1.595 4.925 1.685 ;
        RECT 5.37 1.915 5.46 2.005 ;
        RECT 5.555 1.595 5.645 1.685 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 1.965 3.065 2.065 3.76 ;
        RECT 4.33 3.2 4.43 3.76 ;
        RECT 5 3.23 5.1 3.76 ;
        RECT 5.63 3.065 5.73 3.76 ;
        RECT 0 3.44 5.8 3.76 ;
        RECT 1.65 -0.16 1.75 0.535 ;
        RECT 3.685 -0.16 3.785 0.56 ;
        RECT 4.24 -0.16 4.34 0.56 ;
        RECT 5.125 -0.16 5.225 0.535 ;
        RECT 0 -0.16 5.8 0.16 ;
      LAYER CUT01 ;
        RECT 1.655 0.405 1.745 0.495 ;
        RECT 1.655 0.205 1.745 0.295 ;
        RECT 1.97 3.305 2.06 3.395 ;
        RECT 1.97 3.105 2.06 3.195 ;
        RECT 3.69 0.43 3.78 0.52 ;
        RECT 3.69 0.23 3.78 0.32 ;
        RECT 4.245 0.43 4.335 0.52 ;
        RECT 4.245 0.23 4.335 0.32 ;
        RECT 4.335 3.245 4.425 3.335 ;
        RECT 5.005 3.275 5.095 3.365 ;
        RECT 5.13 0.405 5.22 0.495 ;
        RECT 5.13 0.205 5.22 0.295 ;
        RECT 5.635 3.305 5.725 3.395 ;
        RECT 5.635 3.105 5.725 3.195 ;
    END
  END VSS
  PIN VYY
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT 1.5 0.78 2.5 2.82 ;
      LAYER MET1 ;
        RECT 1.65 2.125 1.75 2.46 ;
        RECT 1.965 2.125 2.065 2.46 ;
        RECT 0.06 2.125 5.74 2.275 ;
        RECT 1.65 1.14 1.75 1.475 ;
        RECT 0.06 1.325 5.74 1.475 ;
      LAYER CUT01 ;
        RECT 1.655 2.33 1.745 2.42 ;
        RECT 1.655 2.13 1.745 2.22 ;
        RECT 1.655 1.38 1.745 1.47 ;
        RECT 1.655 1.18 1.745 1.27 ;
        RECT 1.97 2.33 2.06 2.42 ;
        RECT 1.97 2.13 2.06 2.22 ;
    END
  END VYY
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4477 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 3.91 0.3 4.08 1.185 ;
        RECT 3.91 0.7 4.67 0.9 ;
        RECT 4.5 0.3 4.67 1.185 ;
      LAYER CUT01 ;
        RECT 3.95 1.075 4.04 1.165 ;
        RECT 3.95 0.505 4.04 0.595 ;
        RECT 3.95 0.305 4.04 0.395 ;
        RECT 4.54 1.075 4.63 1.165 ;
        RECT 4.54 0.505 4.63 0.595 ;
        RECT 4.54 0.305 4.63 0.395 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT 0.5 -0.5 1.5 4.1 ;
        RECT 2.5 -0.5 3.5 4.1 ;
        RECT -0.5 -0.5 6.3 0.78 ;
        RECT -0.5 2.82 6.3 4.1 ;
    END
  END VPW
  OBS
    LAYER MET1 ;
      RECT 1.91 0.385 2.36 0.485 ;
      RECT 1.91 0.285 2.01 1.225 ;
      RECT 1.865 1.125 3.575 1.225 ;
      RECT 2.18 2.375 2.37 2.475 ;
      RECT 4.13 2.975 4.7 3.075 ;
      RECT 4.13 2.975 4.23 3.28 ;
      RECT 2.225 3.18 4.23 3.28 ;
      RECT 2.225 2.375 2.325 3.315 ;
      RECT 3.53 2.375 3.825 2.475 ;
      RECT 3.93 2.775 5.145 2.875 ;
      RECT 3.53 2.375 3.63 3.08 ;
      RECT 3.93 2.775 4.03 3.08 ;
      RECT 3.53 2.98 4.03 3.08 ;
      RECT 3.73 2.575 5.47 2.675 ;
      RECT 4.8 3.01 5.47 3.11 ;
      RECT 4.8 3.01 4.9 3.275 ;
      RECT 4.6 3.175 4.9 3.275 ;
      RECT 5.37 2.575 5.47 3.315 ;
      RECT 4.865 0.285 4.965 1.225 ;
      RECT 4.865 1.125 5.48 1.225 ;
      RECT 4.135 2.375 5.73 2.475 ;
      RECT 5.63 2.375 5.73 2.565 ;
  END
END SC22LSBIORCLXL1

MACRO SC22LSBIORCLXP1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSBIORCLXP1 0 0 ;
  SIZE 7.4 BY 3.6 ;
  SYMMETRY X Y ;
  SITE WCORE3600 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.117 LAYER MET1 ;
    ANTENNAMAXCUTCAR 25.643162 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VYY ;
    PORT
      LAYER MET1 ;
        RECT 1.3 0.4 1.4 0.85 ;
        RECT 1.3 0.74 1.81 0.85 ;
      LAYER CUT01 ;
        RECT 1.305 0.45 1.395 0.54 ;
        RECT 1.675 0.745 1.765 0.835 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.0845 LAYER MET1 ;
    ANTENNAMAXCUTCAR 35.505803 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 7 0.4 7.1 0.85 ;
        RECT 6.5 0.75 7.1 0.85 ;
      LAYER CUT01 ;
        RECT 6.545 0.755 6.635 0.845 ;
        RECT 7.005 0.45 7.095 0.54 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 0.5 2.82 ;
        RECT 3.7 0.78 7.9 2.82 ;
      LAYER MET1 ;
        RECT 3.81 1.595 3.99 1.96 ;
        RECT 4.4 1.595 4.58 1.96 ;
        RECT 4.99 1.595 5.17 1.96 ;
        RECT 5.58 1.595 5.76 1.96 ;
        RECT 6.17 1.595 6.35 1.96 ;
        RECT 6.395 1.64 6.575 2.005 ;
        RECT 6.7 1.595 6.88 1.96 ;
        RECT 6.925 1.64 7.105 2.005 ;
        RECT 7.11 1.595 7.29 1.96 ;
        RECT 0 1.64 7.4 1.96 ;
      LAYER CUT01 ;
        RECT 0.175 1.86 0.265 1.95 ;
        RECT 0.175 1.65 0.265 1.74 ;
        RECT 3.855 1.595 3.945 1.685 ;
        RECT 4.445 1.595 4.535 1.685 ;
        RECT 5.035 1.595 5.125 1.685 ;
        RECT 5.625 1.595 5.715 1.685 ;
        RECT 6.215 1.595 6.305 1.685 ;
        RECT 6.44 1.915 6.53 2.005 ;
        RECT 6.745 1.595 6.835 1.685 ;
        RECT 6.97 1.915 7.06 2.005 ;
        RECT 7.155 1.595 7.245 1.685 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 1.93 3.065 2.03 3.76 ;
        RECT 2.45 3.065 2.55 3.76 ;
        RECT 4.51 3.23 4.61 3.76 ;
        RECT 5.045 3.395 5.225 3.76 ;
        RECT 5.375 3.395 5.555 3.76 ;
        RECT 6.07 3.23 6.17 3.76 ;
        RECT 6.44 3.23 6.54 3.76 ;
        RECT 6.96 3.065 7.06 3.76 ;
        RECT 0 3.44 7.4 3.76 ;
        RECT 1.65 -0.16 1.75 0.535 ;
        RECT 2.17 -0.16 2.27 0.535 ;
        RECT 3.885 -0.16 3.985 0.56 ;
        RECT 4.44 -0.16 4.54 0.56 ;
        RECT 5.03 -0.16 5.13 0.56 ;
        RECT 5.585 -0.16 5.685 0.56 ;
        RECT 6.215 -0.16 6.315 0.43 ;
        RECT 6.735 -0.16 6.835 0.43 ;
        RECT 0 -0.16 7.4 0.16 ;
      LAYER CUT01 ;
        RECT 1.655 0.405 1.745 0.495 ;
        RECT 1.655 0.205 1.745 0.295 ;
        RECT 1.935 3.305 2.025 3.395 ;
        RECT 1.935 3.105 2.025 3.195 ;
        RECT 2.175 0.405 2.265 0.495 ;
        RECT 2.175 0.205 2.265 0.295 ;
        RECT 2.455 3.305 2.545 3.395 ;
        RECT 2.455 3.105 2.545 3.195 ;
        RECT 3.89 0.43 3.98 0.52 ;
        RECT 3.89 0.23 3.98 0.32 ;
        RECT 4.445 0.43 4.535 0.52 ;
        RECT 4.445 0.23 4.535 0.32 ;
        RECT 4.515 3.275 4.605 3.365 ;
        RECT 5.035 0.43 5.125 0.52 ;
        RECT 5.035 0.23 5.125 0.32 ;
        RECT 5.09 3.395 5.18 3.485 ;
        RECT 5.42 3.395 5.51 3.485 ;
        RECT 5.59 0.43 5.68 0.52 ;
        RECT 5.59 0.23 5.68 0.32 ;
        RECT 6.075 3.275 6.165 3.365 ;
        RECT 6.22 0.295 6.31 0.385 ;
        RECT 6.445 3.275 6.535 3.365 ;
        RECT 6.74 0.295 6.83 0.385 ;
        RECT 6.965 3.305 7.055 3.395 ;
        RECT 6.965 3.105 7.055 3.195 ;
    END
  END VSS
  PIN VYY
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT 1.5 0.78 2.7 2.82 ;
      LAYER MET1 ;
        RECT 1.65 2.125 1.75 2.46 ;
        RECT 1.93 2.125 2.03 2.46 ;
        RECT 2.45 2.125 2.55 2.46 ;
        RECT 0.06 2.125 7.34 2.275 ;
        RECT 1.65 1.14 1.75 1.475 ;
        RECT 2.17 1.14 2.27 1.475 ;
        RECT 0.06 1.325 7.34 1.475 ;
      LAYER CUT01 ;
        RECT 1.655 2.33 1.745 2.42 ;
        RECT 1.655 2.13 1.745 2.22 ;
        RECT 1.655 1.38 1.745 1.47 ;
        RECT 1.655 1.18 1.745 1.27 ;
        RECT 1.935 2.33 2.025 2.42 ;
        RECT 1.935 2.13 2.025 2.22 ;
        RECT 2.175 1.38 2.265 1.47 ;
        RECT 2.175 1.18 2.265 1.27 ;
        RECT 2.455 2.33 2.545 2.42 ;
        RECT 2.455 2.13 2.545 2.22 ;
    END
  END VYY
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.824 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 4.11 0.3 4.28 1.185 ;
        RECT 4.7 0.3 4.87 1.185 ;
        RECT 5.29 0.3 5.46 1.185 ;
        RECT 4.11 0.75 6.05 1.05 ;
        RECT 5.88 0.75 6.05 1.185 ;
      LAYER CUT01 ;
        RECT 4.15 1.075 4.24 1.165 ;
        RECT 4.15 0.505 4.24 0.595 ;
        RECT 4.15 0.305 4.24 0.395 ;
        RECT 4.74 1.075 4.83 1.165 ;
        RECT 4.74 0.505 4.83 0.595 ;
        RECT 4.74 0.305 4.83 0.395 ;
        RECT 5.33 1.075 5.42 1.165 ;
        RECT 5.33 0.505 5.42 0.595 ;
        RECT 5.33 0.305 5.42 0.395 ;
        RECT 5.92 1.075 6.01 1.165 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT 0.5 -0.5 1.5 4.1 ;
        RECT 2.7 -0.5 3.7 4.1 ;
        RECT -0.5 -0.5 7.9 0.78 ;
        RECT -0.5 2.82 7.9 4.1 ;
    END
  END VPW
  OBS
    LAYER MET1 ;
      RECT 1.91 0.785 2.63 0.885 ;
      RECT 1.91 0.285 2.01 1.225 ;
      RECT 2.53 0.4 2.63 1.225 ;
      RECT 1.865 1.125 2.055 1.225 ;
      RECT 2.53 1.125 2.815 1.225 ;
      RECT 2.145 2.375 2.335 2.475 ;
      RECT 2.19 2.8 2.87 2.9 ;
      RECT 4.31 2.975 5.77 3.075 ;
      RECT 2.77 2.8 2.87 3.28 ;
      RECT 4.31 2.975 4.41 3.28 ;
      RECT 2.77 3.18 4.41 3.28 ;
      RECT 2.19 2.375 2.29 3.315 ;
      RECT 3.44 2.375 4.005 2.475 ;
      RECT 4.11 2.775 6.215 2.875 ;
      RECT 3.44 2.375 3.54 3.08 ;
      RECT 4.11 2.775 4.21 3.08 ;
      RECT 3.44 2.98 4.21 3.08 ;
      RECT 3.64 2.575 6.8 2.675 ;
      RECT 3.64 2.575 3.825 2.685 ;
      RECT 5.87 3 6.8 3.1 ;
      RECT 5.87 3 5.97 3.275 ;
      RECT 4.75 3.175 5.97 3.275 ;
      RECT 6.7 2.575 6.8 3.315 ;
      RECT 6.475 0.4 6.575 0.64 ;
      RECT 6.3 0.54 6.575 0.64 ;
      RECT 6.3 0.54 6.4 1.225 ;
      RECT 6.3 1.125 7.08 1.225 ;
      RECT 4.285 2.375 7.33 2.475 ;
      RECT 7.23 2.375 7.33 2.565 ;
  END
END SC22LSBIORCLXP1

MACRO SC22LSBOANDCLXL1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSBOANDCLXL1 0 0 ;
  SIZE 5.6 BY 3.6 ;
  SYMMETRY X Y ;
  SITE WCORE3600 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.0585 LAYER MET1 ;
    ANTENNAMAXCUTCAR 51.286325 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.62 0.4 0.72 0.85 ;
        RECT 0.3 0.74 0.72 0.85 ;
      LAYER CUT01 ;
        RECT 0.345 0.745 0.435 0.835 ;
        RECT 0.625 0.45 0.715 0.54 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.0585 LAYER MET1 ;
    ANTENNAMAXCUTCAR 51.286325 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VYY ;
    PORT
      LAYER MET1 ;
        RECT 3.55 0.4 3.65 1.225 ;
        RECT 3.55 1.125 3.88 1.225 ;
      LAYER CUT01 ;
        RECT 3.555 0.45 3.645 0.54 ;
        RECT 3.745 1.13 3.835 1.22 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 0.94 2.82 ;
        RECT 5.1 0.78 6.1 2.82 ;
      LAYER MET1 ;
        RECT 0.095 1.64 0.275 2.005 ;
        RECT 0.325 1.595 0.505 1.96 ;
        RECT 0.65 1.64 0.83 2.005 ;
        RECT 0 1.64 5.6 1.96 ;
      LAYER CUT01 ;
        RECT 0.14 1.915 0.23 2.005 ;
        RECT 0.37 1.595 0.46 1.685 ;
        RECT 0.695 1.915 0.785 2.005 ;
        RECT 5.335 1.86 5.425 1.95 ;
        RECT 5.335 1.65 5.425 1.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.685 3.065 0.785 3.76 ;
        RECT 3.84 3.245 3.94 3.76 ;
        RECT 0 3.44 5.6 3.76 ;
        RECT 0.36 -0.16 0.46 0.535 ;
        RECT 2.115 -0.16 2.215 0.56 ;
        RECT 2.65 -0.16 2.75 0.56 ;
        RECT 0 -0.16 5.6 0.16 ;
      LAYER CUT01 ;
        RECT 0.365 0.405 0.455 0.495 ;
        RECT 0.365 0.205 0.455 0.295 ;
        RECT 0.69 3.305 0.78 3.395 ;
        RECT 0.69 3.105 0.78 3.195 ;
        RECT 2.12 0.43 2.21 0.52 ;
        RECT 2.12 0.23 2.21 0.32 ;
        RECT 2.655 0.43 2.745 0.52 ;
        RECT 2.655 0.23 2.745 0.32 ;
        RECT 3.845 3.295 3.935 3.385 ;
    END
  END VSS
  PIN VYY
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT 1.94 0.78 4.1 2.82 ;
      LAYER MET1 ;
        RECT 0.06 2.125 5.54 2.275 ;
        RECT 2.115 1.14 2.215 1.475 ;
        RECT 2.65 1.14 2.75 1.475 ;
        RECT 3.185 1.14 3.285 1.475 ;
        RECT 0.06 1.325 5.54 1.475 ;
      LAYER CUT01 ;
        RECT 2.12 1.38 2.21 1.47 ;
        RECT 2.12 1.18 2.21 1.27 ;
        RECT 2.65 2.155 2.74 2.245 ;
        RECT 2.655 1.38 2.745 1.47 ;
        RECT 2.655 1.18 2.745 1.27 ;
        RECT 3.19 1.38 3.28 1.47 ;
        RECT 3.19 1.18 3.28 1.27 ;
        RECT 3.535 1.355 3.625 1.445 ;
        RECT 3.575 2.155 3.665 2.245 ;
    END
  END VYY
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4477 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 2.34 0.3 2.51 1.185 ;
        RECT 2.34 0.7 3.06 0.9 ;
        RECT 2.89 0.3 3.06 1.185 ;
      LAYER CUT01 ;
        RECT 2.38 1.075 2.47 1.165 ;
        RECT 2.38 0.505 2.47 0.595 ;
        RECT 2.38 0.305 2.47 0.395 ;
        RECT 2.93 1.075 3.02 1.165 ;
        RECT 2.93 0.505 3.02 0.595 ;
        RECT 2.93 0.305 3.02 0.395 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT 0.94 -0.5 1.94 4.1 ;
        RECT 4.1 -0.5 5.1 4.1 ;
        RECT -0.5 -0.5 6.1 0.78 ;
        RECT -0.5 2.82 6.1 4.1 ;
    END
  END VPW
  OBS
    LAYER MET1 ;
      RECT 0.1 0.285 0.2 1.225 ;
      RECT 0.86 0.4 0.96 1.225 ;
      RECT 0.06 1.125 2.015 1.225 ;
      RECT 2.98 2.77 3.245 2.87 ;
      RECT 0.425 2.8 1.11 2.9 ;
      RECT 2.98 2.77 3.08 3.075 ;
      RECT 2.495 2.975 3.08 3.075 ;
      RECT 1.01 2.8 1.11 3.28 ;
      RECT 2.495 2.975 2.595 3.28 ;
      RECT 1.01 3.18 2.595 3.28 ;
      RECT 0.425 2.415 0.525 3.315 ;
      RECT 1.96 2.375 2.255 2.475 ;
      RECT 2.77 2.575 3.5 2.675 ;
      RECT 3.4 2.575 3.5 2.87 ;
      RECT 3.4 2.77 3.61 2.87 ;
      RECT 2.77 2.575 2.87 2.875 ;
      RECT 2.295 2.775 2.87 2.875 ;
      RECT 1.96 2.375 2.06 3.085 ;
      RECT 2.295 2.775 2.395 3.085 ;
      RECT 1.96 2.985 2.395 3.085 ;
      RECT 2.695 3.19 3.72 3.29 ;
      RECT 2.445 2.375 3.94 2.475 ;
      RECT 2.445 2.375 2.545 2.675 ;
      RECT 2.16 2.575 2.545 2.675 ;
      RECT 3.84 2.375 3.94 3.09 ;
      RECT 3.195 2.99 3.94 3.09 ;
  END
END SC22LSBOANDCLXL1

MACRO SC22LSBOANDCLXP1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSBOANDCLXP1 0 0 ;
  SIZE 7.2 BY 3.6 ;
  SYMMETRY X Y ;
  SITE WCORE3600 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.117 LAYER MET1 ;
    ANTENNAMAXCUTCAR 25.643162 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 1 0.4 1.1 0.85 ;
        RECT 0.58 0.74 1.1 0.85 ;
      LAYER CUT01 ;
        RECT 0.625 0.745 0.715 0.835 ;
        RECT 1.005 0.45 1.095 0.54 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.117 LAYER MET1 ;
    ANTENNAMAXCUTCAR 32.00256 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VYY ;
    PORT
      LAYER MET1 ;
        RECT 5.15 0.4 5.25 1.225 ;
        RECT 5.105 1.125 5.295 1.225 ;
      LAYER CUT01 ;
        RECT 5.155 1.13 5.245 1.22 ;
        RECT 5.155 0.45 5.245 0.54 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 1.245 2.82 ;
        RECT 6.7 0.78 7.7 2.82 ;
      LAYER MET1 ;
        RECT 0.075 1.595 0.255 1.96 ;
        RECT 0.095 1.64 0.275 2.005 ;
        RECT 0.395 1.64 0.575 2.005 ;
        RECT 0.635 1.595 0.815 1.96 ;
        RECT 0.955 1.64 1.135 2.005 ;
        RECT 0 1.64 7.2 1.96 ;
      LAYER CUT01 ;
        RECT 0.12 1.595 0.21 1.685 ;
        RECT 0.14 1.915 0.23 2.005 ;
        RECT 0.44 1.915 0.53 2.005 ;
        RECT 0.68 1.595 0.77 1.685 ;
        RECT 1 1.915 1.09 2.005 ;
        RECT 6.935 1.86 7.025 1.95 ;
        RECT 6.935 1.65 7.025 1.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.47 3.065 0.57 3.76 ;
        RECT 0.99 3.065 1.09 3.76 ;
        RECT 4.795 3.41 4.975 3.76 ;
        RECT 5.39 3.065 5.49 3.76 ;
        RECT 0 3.44 7.2 3.76 ;
        RECT 0.12 -0.16 0.22 0.535 ;
        RECT 0.64 -0.16 0.74 0.535 ;
        RECT 2.405 -0.16 2.505 0.56 ;
        RECT 2.94 -0.16 3.04 0.56 ;
        RECT 3.49 -0.16 3.59 0.56 ;
        RECT 4.025 -0.16 4.125 0.56 ;
        RECT 0 -0.16 7.2 0.16 ;
      LAYER CUT01 ;
        RECT 0.125 0.405 0.215 0.495 ;
        RECT 0.125 0.205 0.215 0.295 ;
        RECT 0.475 3.305 0.565 3.395 ;
        RECT 0.475 3.105 0.565 3.195 ;
        RECT 0.645 0.405 0.735 0.495 ;
        RECT 0.645 0.205 0.735 0.295 ;
        RECT 0.995 3.305 1.085 3.395 ;
        RECT 0.995 3.105 1.085 3.195 ;
        RECT 2.41 0.43 2.5 0.52 ;
        RECT 2.41 0.23 2.5 0.32 ;
        RECT 2.945 0.43 3.035 0.52 ;
        RECT 2.945 0.23 3.035 0.32 ;
        RECT 3.495 0.43 3.585 0.52 ;
        RECT 3.495 0.23 3.585 0.32 ;
        RECT 4.03 0.43 4.12 0.52 ;
        RECT 4.03 0.23 4.12 0.32 ;
        RECT 4.84 3.41 4.93 3.5 ;
        RECT 5.395 3.305 5.485 3.395 ;
        RECT 5.395 3.105 5.485 3.195 ;
    END
  END VSS
  PIN VYY
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT 2.245 0.78 5.7 2.82 ;
      LAYER MET1 ;
        RECT 5.39 2.125 5.49 2.46 ;
        RECT 0.06 2.125 7.14 2.275 ;
        RECT 2.405 1.14 2.505 1.475 ;
        RECT 4.545 1.14 4.645 1.475 ;
        RECT 4.865 1.14 4.965 1.475 ;
        RECT 0.06 1.325 7.14 1.475 ;
      LAYER CUT01 ;
        RECT 2.41 1.38 2.5 1.47 ;
        RECT 2.41 1.18 2.5 1.27 ;
        RECT 2.945 1.355 3.035 1.445 ;
        RECT 2.965 2.155 3.055 2.245 ;
        RECT 3.495 1.355 3.585 1.445 ;
        RECT 3.885 2.155 3.975 2.245 ;
        RECT 4.03 1.355 4.12 1.445 ;
        RECT 4.55 1.38 4.64 1.47 ;
        RECT 4.55 1.18 4.64 1.27 ;
        RECT 4.84 2.155 4.93 2.245 ;
        RECT 4.87 1.38 4.96 1.47 ;
        RECT 4.87 1.18 4.96 1.27 ;
        RECT 5.395 2.33 5.485 2.42 ;
        RECT 5.395 2.13 5.485 2.22 ;
    END
  END VYY
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.824 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 2.63 0.3 2.8 1.185 ;
        RECT 3.18 0.3 3.35 1.185 ;
        RECT 3.73 0.3 3.9 1.185 ;
        RECT 2.63 0.75 4.42 1.05 ;
        RECT 4.25 0.75 4.42 1.185 ;
      LAYER CUT01 ;
        RECT 2.67 1.075 2.76 1.165 ;
        RECT 2.67 0.505 2.76 0.595 ;
        RECT 2.67 0.305 2.76 0.395 ;
        RECT 3.22 1.075 3.31 1.165 ;
        RECT 3.22 0.505 3.31 0.595 ;
        RECT 3.22 0.305 3.31 0.395 ;
        RECT 3.77 1.075 3.86 1.165 ;
        RECT 3.77 0.505 3.86 0.595 ;
        RECT 3.77 0.305 3.86 0.395 ;
        RECT 4.29 1.075 4.38 1.165 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT 1.245 -0.5 2.245 4.1 ;
        RECT 5.7 -0.5 6.7 4.1 ;
        RECT -0.5 -0.5 7.7 0.78 ;
        RECT -0.5 2.82 7.7 4.1 ;
    END
  END VPW
  OBS
    LAYER MET1 ;
      RECT 0.38 0.285 0.48 1.225 ;
      RECT 1.26 0.4 1.36 1.225 ;
      RECT 0.335 1.125 1.36 1.225 ;
      RECT 0.685 2.375 0.875 2.475 ;
      RECT 3.38 2.775 3.56 2.875 ;
      RECT 4.1 2.775 4.485 2.875 ;
      RECT 0.73 2.8 1.415 2.9 ;
      RECT 3.42 2.775 3.52 3.075 ;
      RECT 4.1 2.775 4.2 3.075 ;
      RECT 2.875 2.975 4.2 3.075 ;
      RECT 1.315 2.8 1.415 3.28 ;
      RECT 2.875 2.975 2.975 3.28 ;
      RECT 1.315 3.18 2.975 3.28 ;
      RECT 0.73 2.375 0.83 3.315 ;
      RECT 1.995 2.375 2.57 2.475 ;
      RECT 3.095 2.575 4.82 2.675 ;
      RECT 3.86 2.575 3.96 2.875 ;
      RECT 3.095 2.575 3.195 2.875 ;
      RECT 2.675 2.775 3.195 2.875 ;
      RECT 3.82 2.775 4 2.875 ;
      RECT 4.72 2.575 4.82 2.89 ;
      RECT 1.995 2.375 2.095 3.08 ;
      RECT 2.675 2.775 2.775 3.08 ;
      RECT 1.995 2.98 2.775 3.08 ;
      RECT 2.76 2.375 5.23 2.475 ;
      RECT 2.76 2.375 2.86 2.675 ;
      RECT 2.195 2.575 2.86 2.675 ;
      RECT 5.13 2.375 5.23 3.09 ;
      RECT 4.3 2.99 5.23 3.09 ;
      RECT 3.075 3.19 5.27 3.29 ;
  END
END SC22LSBOANDCLXP1

MACRO SC22LSBOCLXL1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSBOCLXL1 0 0 ;
  SIZE 5.4 BY 3.6 ;
  SYMMETRY X Y ;
  SITE WCORE3600 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.0585 LAYER MET1 ;
    ANTENNAMAXCUTCAR 51.286325 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.62 0.4 0.72 0.85 ;
        RECT 0.3 0.74 0.72 0.85 ;
      LAYER CUT01 ;
        RECT 0.345 0.745 0.435 0.835 ;
        RECT 0.625 0.45 0.715 0.54 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 0.94 2.82 ;
        RECT 4.9 0.78 5.9 2.82 ;
      LAYER MET1 ;
        RECT 0.095 1.64 0.275 2.005 ;
        RECT 0.325 1.595 0.505 1.96 ;
        RECT 0.65 1.64 0.83 2.005 ;
        RECT 0 1.64 5.4 1.96 ;
      LAYER CUT01 ;
        RECT 0.14 1.915 0.23 2.005 ;
        RECT 0.37 1.595 0.46 1.685 ;
        RECT 0.695 1.915 0.785 2.005 ;
        RECT 5.135 1.86 5.225 1.95 ;
        RECT 5.135 1.65 5.225 1.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.685 3.065 0.785 3.76 ;
        RECT 2.79 3.2 2.89 3.76 ;
        RECT 0 3.44 5.4 3.76 ;
        RECT 0.36 -0.16 0.46 0.535 ;
        RECT 2.125 -0.16 2.225 0.56 ;
        RECT 2.66 -0.16 2.76 0.56 ;
        RECT 0 -0.16 5.4 0.16 ;
      LAYER CUT01 ;
        RECT 0.365 0.405 0.455 0.495 ;
        RECT 0.365 0.205 0.455 0.295 ;
        RECT 0.69 3.305 0.78 3.395 ;
        RECT 0.69 3.105 0.78 3.195 ;
        RECT 2.13 0.43 2.22 0.52 ;
        RECT 2.13 0.23 2.22 0.32 ;
        RECT 2.665 0.43 2.755 0.52 ;
        RECT 2.665 0.23 2.755 0.32 ;
        RECT 2.795 3.245 2.885 3.335 ;
    END
  END VSS
  PIN VYY
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT 1.94 0.78 3.9 2.82 ;
      LAYER MET1 ;
        RECT 0.06 2.125 5.34 2.275 ;
        RECT 2.125 1.14 2.225 1.475 ;
        RECT 2.66 1.14 2.76 1.475 ;
        RECT 3.195 1.14 3.295 1.475 ;
        RECT 3.65 1.14 3.75 1.475 ;
        RECT 0.06 1.325 5.34 1.475 ;
      LAYER CUT01 ;
        RECT 2.13 1.38 2.22 1.47 ;
        RECT 2.13 1.18 2.22 1.27 ;
        RECT 2.635 2.155 2.725 2.245 ;
        RECT 2.665 1.38 2.755 1.47 ;
        RECT 2.665 1.18 2.755 1.27 ;
        RECT 3.2 1.38 3.29 1.47 ;
        RECT 3.2 1.18 3.29 1.27 ;
        RECT 3.555 2.155 3.645 2.245 ;
        RECT 3.655 1.38 3.745 1.47 ;
        RECT 3.655 1.18 3.745 1.27 ;
    END
  END VYY
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4477 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 2.35 0.3 2.52 1.185 ;
        RECT 2.35 0.7 3.07 0.9 ;
        RECT 2.9 0.3 3.07 1.185 ;
      LAYER CUT01 ;
        RECT 2.39 1.075 2.48 1.165 ;
        RECT 2.39 0.505 2.48 0.595 ;
        RECT 2.39 0.305 2.48 0.395 ;
        RECT 2.94 1.075 3.03 1.165 ;
        RECT 2.94 0.505 3.03 0.595 ;
        RECT 2.94 0.305 3.03 0.395 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT 0.94 -0.5 1.94 4.1 ;
        RECT 3.9 -0.5 4.9 4.1 ;
        RECT -0.5 -0.5 5.9 0.78 ;
        RECT -0.5 2.82 5.9 4.1 ;
    END
  END VPW
  OBS
    LAYER MET1 ;
      RECT 0.1 0.285 0.2 1.225 ;
      RECT 0.86 0.4 0.96 1.225 ;
      RECT 0.06 1.125 2.025 1.225 ;
      RECT 2.985 2.77 3.215 2.87 ;
      RECT 0.425 2.8 1.11 2.9 ;
      RECT 2.985 2.77 3.085 3.075 ;
      RECT 2.58 2.975 3.085 3.075 ;
      RECT 1.01 2.8 1.11 3.28 ;
      RECT 2.58 2.975 2.68 3.28 ;
      RECT 1.01 3.18 2.68 3.28 ;
      RECT 0.425 2.415 0.525 3.315 ;
      RECT 1.97 2.375 2.265 2.475 ;
      RECT 2.765 2.575 3.55 2.675 ;
      RECT 2.765 2.575 2.865 2.875 ;
      RECT 2.37 2.775 2.865 2.875 ;
      RECT 3.45 2.575 3.55 2.925 ;
      RECT 1.97 2.375 2.07 3.08 ;
      RECT 2.37 2.775 2.47 3.08 ;
      RECT 1.97 2.98 2.47 3.08 ;
      RECT 2.455 2.375 3.75 2.475 ;
      RECT 2.455 2.375 2.555 2.675 ;
      RECT 2.17 2.575 2.555 2.675 ;
      RECT 3.65 2.375 3.75 3.275 ;
      RECT 3.05 3.175 3.75 3.275 ;
  END
END SC22LSBOCLXL1

MACRO SC22LSBOCLXP1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSBOCLXP1 0 0 ;
  SIZE 6.6 BY 3.6 ;
  SYMMETRY X Y ;
  SITE WCORE3600 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.117 LAYER MET1 ;
    ANTENNAMAXCUTCAR 25.643162 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 1 0.4 1.1 0.85 ;
        RECT 0.58 0.74 1.1 0.85 ;
      LAYER CUT01 ;
        RECT 0.625 0.745 0.715 0.835 ;
        RECT 1.005 0.45 1.095 0.54 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 1.245 2.82 ;
        RECT 6.1 0.78 7.1 2.82 ;
      LAYER MET1 ;
        RECT 0.075 1.595 0.255 1.96 ;
        RECT 0.095 1.64 0.275 2.005 ;
        RECT 0.395 1.64 0.575 2.005 ;
        RECT 0.635 1.595 0.815 1.96 ;
        RECT 0.955 1.64 1.135 2.005 ;
        RECT 0 1.64 6.6 1.96 ;
      LAYER CUT01 ;
        RECT 0.12 1.595 0.21 1.685 ;
        RECT 0.14 1.915 0.23 2.005 ;
        RECT 0.44 1.915 0.53 2.005 ;
        RECT 0.68 1.595 0.77 1.685 ;
        RECT 1 1.915 1.09 2.005 ;
        RECT 6.335 1.86 6.425 1.95 ;
        RECT 6.335 1.65 6.425 1.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.47 3.065 0.57 3.76 ;
        RECT 0.99 3.065 1.09 3.76 ;
        RECT 3.075 3.25 3.175 3.76 ;
        RECT 4.055 3.25 4.155 3.76 ;
        RECT 4.575 3.25 4.675 3.76 ;
        RECT 0 3.44 6.6 3.76 ;
        RECT 0.12 -0.16 0.22 0.535 ;
        RECT 0.64 -0.16 0.74 0.535 ;
        RECT 2.395 -0.16 2.495 0.56 ;
        RECT 2.93 -0.16 3.03 0.56 ;
        RECT 3.48 -0.16 3.58 0.56 ;
        RECT 4.015 -0.16 4.115 0.56 ;
        RECT 0 -0.16 6.6 0.16 ;
      LAYER CUT01 ;
        RECT 0.125 0.405 0.215 0.495 ;
        RECT 0.125 0.205 0.215 0.295 ;
        RECT 0.475 3.305 0.565 3.395 ;
        RECT 0.475 3.105 0.565 3.195 ;
        RECT 0.645 0.405 0.735 0.495 ;
        RECT 0.645 0.205 0.735 0.295 ;
        RECT 0.995 3.305 1.085 3.395 ;
        RECT 0.995 3.105 1.085 3.195 ;
        RECT 2.4 0.43 2.49 0.52 ;
        RECT 2.4 0.23 2.49 0.32 ;
        RECT 2.935 0.43 3.025 0.52 ;
        RECT 2.935 0.23 3.025 0.32 ;
        RECT 3.08 3.295 3.17 3.385 ;
        RECT 3.485 0.43 3.575 0.52 ;
        RECT 3.485 0.23 3.575 0.32 ;
        RECT 4.02 0.43 4.11 0.52 ;
        RECT 4.02 0.23 4.11 0.32 ;
        RECT 4.06 3.295 4.15 3.385 ;
        RECT 4.58 3.295 4.67 3.385 ;
    END
  END VSS
  PIN VYY
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT 2.245 0.78 5.1 2.82 ;
      LAYER MET1 ;
        RECT 0.06 2.125 6.54 2.275 ;
        RECT 2.395 1.14 2.495 1.475 ;
        RECT 4.535 1.14 4.635 1.475 ;
        RECT 4.85 1.14 4.95 1.475 ;
        RECT 0.06 1.325 6.54 1.475 ;
      LAYER CUT01 ;
        RECT 2.4 1.38 2.49 1.47 ;
        RECT 2.4 1.18 2.49 1.27 ;
        RECT 2.935 1.355 3.025 1.445 ;
        RECT 2.94 2.155 3.03 2.245 ;
        RECT 3.485 1.355 3.575 1.445 ;
        RECT 3.86 2.155 3.95 2.245 ;
        RECT 4.02 1.355 4.11 1.445 ;
        RECT 4.54 1.38 4.63 1.47 ;
        RECT 4.54 1.18 4.63 1.27 ;
        RECT 4.78 2.155 4.87 2.245 ;
        RECT 4.855 1.38 4.945 1.47 ;
        RECT 4.855 1.18 4.945 1.27 ;
    END
  END VYY
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.824 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 2.62 0.3 2.79 1.185 ;
        RECT 3.17 0.3 3.34 1.185 ;
        RECT 3.72 0.3 3.89 1.185 ;
        RECT 2.62 0.75 4.41 1.05 ;
        RECT 4.24 0.75 4.41 1.185 ;
      LAYER CUT01 ;
        RECT 2.66 1.075 2.75 1.165 ;
        RECT 2.66 0.505 2.75 0.595 ;
        RECT 2.66 0.305 2.75 0.395 ;
        RECT 3.21 1.075 3.3 1.165 ;
        RECT 3.21 0.505 3.3 0.595 ;
        RECT 3.21 0.305 3.3 0.395 ;
        RECT 3.76 1.075 3.85 1.165 ;
        RECT 3.76 0.505 3.85 0.595 ;
        RECT 3.76 0.305 3.85 0.395 ;
        RECT 4.28 1.075 4.37 1.165 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT 1.245 -0.5 2.245 4.1 ;
        RECT 5.1 -0.5 6.1 4.1 ;
        RECT -0.5 -0.5 7.1 0.78 ;
        RECT -0.5 2.82 7.1 4.1 ;
    END
  END VPW
  OBS
    LAYER MET1 ;
      RECT 0.38 0.285 0.48 1.225 ;
      RECT 1.26 0.4 1.36 1.225 ;
      RECT 0.335 1.125 1.36 1.225 ;
      RECT 0.685 2.375 0.875 2.475 ;
      RECT 3.355 2.775 3.535 2.875 ;
      RECT 4.075 2.775 4.46 2.875 ;
      RECT 0.73 2.8 1.415 2.9 ;
      RECT 3.395 2.775 3.495 3.075 ;
      RECT 4.075 2.775 4.175 3.075 ;
      RECT 2.875 2.975 4.175 3.075 ;
      RECT 1.315 2.8 1.415 3.28 ;
      RECT 2.875 2.975 2.975 3.28 ;
      RECT 1.315 3.18 2.975 3.28 ;
      RECT 0.73 2.375 0.83 3.315 ;
      RECT 1.985 2.375 2.57 2.475 ;
      RECT 3.07 2.575 4.775 2.675 ;
      RECT 3.835 2.575 3.935 2.875 ;
      RECT 3.07 2.575 3.17 2.875 ;
      RECT 2.675 2.775 3.17 2.875 ;
      RECT 3.795 2.775 3.975 2.875 ;
      RECT 4.675 2.575 4.775 2.91 ;
      RECT 1.985 2.375 2.085 3.08 ;
      RECT 2.675 2.775 2.775 3.08 ;
      RECT 1.985 2.98 2.775 3.08 ;
      RECT 2.76 2.375 4.975 2.475 ;
      RECT 2.76 2.375 2.86 2.675 ;
      RECT 2.185 2.575 2.86 2.675 ;
      RECT 4.875 2.375 4.975 3.13 ;
      RECT 4.275 3.03 4.975 3.13 ;
  END
END SC22LSBOCLXP1

MACRO SC22LSBOORCLXL1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSBOORCLXL1 0 0 ;
  SIZE 5.8 BY 3.6 ;
  SYMMETRY X Y ;
  SITE WCORE3600 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.0585 LAYER MET1 ;
    ANTENNAMAXCUTCAR 51.286325 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.62 0.4 0.72 0.85 ;
        RECT 0.3 0.74 0.72 0.85 ;
      LAYER CUT01 ;
        RECT 0.345 0.745 0.435 0.835 ;
        RECT 0.625 0.45 0.715 0.54 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.0585 LAYER MET1 ;
    ANTENNAMAXCUTCAR 51.286325 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VYY ;
    PORT
      LAYER MET1 ;
        RECT 3.84 0.4 3.94 0.85 ;
        RECT 3.5 0.74 3.94 0.85 ;
      LAYER CUT01 ;
        RECT 3.545 0.745 3.635 0.835 ;
        RECT 3.845 0.45 3.935 0.54 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 0.94 2.82 ;
        RECT 5.3 0.78 6.3 2.82 ;
      LAYER MET1 ;
        RECT 0.095 1.64 0.275 2.005 ;
        RECT 0.325 1.595 0.505 1.96 ;
        RECT 0.65 1.64 0.83 2.005 ;
        RECT 0 1.64 5.8 1.96 ;
      LAYER CUT01 ;
        RECT 0.14 1.915 0.23 2.005 ;
        RECT 0.37 1.595 0.46 1.685 ;
        RECT 0.695 1.915 0.785 2.005 ;
        RECT 5.535 1.86 5.625 1.95 ;
        RECT 5.535 1.65 5.625 1.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.685 3.065 0.785 3.76 ;
        RECT 2.76 3.2 2.86 3.76 ;
        RECT 3.43 3.23 3.53 3.76 ;
        RECT 4.05 3.065 4.15 3.76 ;
        RECT 0 3.44 5.8 3.76 ;
        RECT 0.36 -0.16 0.46 0.535 ;
        RECT 2.115 -0.16 2.215 0.56 ;
        RECT 2.65 -0.16 2.75 0.56 ;
        RECT 3.56 -0.16 3.66 0.535 ;
        RECT 0 -0.16 5.8 0.16 ;
      LAYER CUT01 ;
        RECT 0.365 0.405 0.455 0.495 ;
        RECT 0.365 0.205 0.455 0.295 ;
        RECT 0.69 3.305 0.78 3.395 ;
        RECT 0.69 3.105 0.78 3.195 ;
        RECT 2.12 0.43 2.21 0.52 ;
        RECT 2.12 0.23 2.21 0.32 ;
        RECT 2.655 0.43 2.745 0.52 ;
        RECT 2.655 0.23 2.745 0.32 ;
        RECT 2.765 3.245 2.855 3.335 ;
        RECT 3.435 3.275 3.525 3.365 ;
        RECT 3.565 0.405 3.655 0.495 ;
        RECT 3.565 0.205 3.655 0.295 ;
        RECT 4.055 3.305 4.145 3.395 ;
        RECT 4.055 3.105 4.145 3.195 ;
    END
  END VSS
  PIN VYY
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT 1.94 0.78 4.3 2.82 ;
      LAYER MET1 ;
        RECT 0.06 2.125 5.74 2.275 ;
        RECT 2.115 1.14 2.215 1.475 ;
        RECT 2.65 1.14 2.75 1.475 ;
        RECT 3.2 1.145 3.3 1.475 ;
        RECT 4.05 1.14 4.15 1.475 ;
        RECT 0.06 1.325 5.74 1.475 ;
      LAYER CUT01 ;
        RECT 2.12 1.38 2.21 1.47 ;
        RECT 2.12 1.18 2.21 1.27 ;
        RECT 2.655 1.38 2.745 1.47 ;
        RECT 2.655 1.18 2.745 1.27 ;
        RECT 3.205 1.385 3.295 1.475 ;
        RECT 3.205 1.185 3.295 1.275 ;
        RECT 3.795 2.155 3.885 2.245 ;
        RECT 4.055 1.38 4.145 1.47 ;
        RECT 4.055 1.18 4.145 1.27 ;
    END
  END VYY
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4477 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 2.34 0.3 2.51 1.185 ;
        RECT 2.34 0.7 3.06 0.9 ;
        RECT 2.89 0.3 3.06 1.185 ;
      LAYER CUT01 ;
        RECT 2.38 1.075 2.47 1.165 ;
        RECT 2.38 0.505 2.47 0.595 ;
        RECT 2.38 0.305 2.47 0.395 ;
        RECT 2.93 1.075 3.02 1.165 ;
        RECT 2.93 0.505 3.02 0.595 ;
        RECT 2.93 0.305 3.02 0.395 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT 0.94 -0.5 1.94 4.1 ;
        RECT 4.3 -0.5 5.3 4.1 ;
        RECT -0.5 -0.5 6.3 0.78 ;
        RECT -0.5 2.82 6.3 4.1 ;
    END
  END VPW
  OBS
    LAYER MET1 ;
      RECT 0.1 0.285 0.2 1.225 ;
      RECT 0.86 0.4 0.96 1.225 ;
      RECT 0.06 1.125 2.015 1.225 ;
      RECT 0.425 2.8 1.11 2.9 ;
      RECT 2.56 2.975 3.13 3.075 ;
      RECT 1.01 2.8 1.11 3.28 ;
      RECT 2.56 2.975 2.66 3.28 ;
      RECT 1.01 3.18 2.66 3.28 ;
      RECT 0.425 2.415 0.525 3.315 ;
      RECT 1.96 2.375 2.255 2.475 ;
      RECT 2.36 2.775 3.575 2.875 ;
      RECT 1.96 2.375 2.06 3.08 ;
      RECT 2.36 2.775 2.46 3.08 ;
      RECT 1.96 2.98 2.46 3.08 ;
      RECT 2.16 2.575 3.89 2.675 ;
      RECT 3.23 3.01 3.89 3.11 ;
      RECT 3.23 3.01 3.33 3.275 ;
      RECT 3.03 3.175 3.33 3.275 ;
      RECT 3.79 2.575 3.89 3.315 ;
      RECT 3.3 0.285 3.4 1.05 ;
      RECT 3.3 0.95 3.66 1.05 ;
      RECT 3.56 0.95 3.66 1.225 ;
      RECT 3.56 1.125 3.925 1.225 ;
      RECT 2.565 2.375 4.195 2.475 ;
  END
END SC22LSBOORCLXL1

MACRO SC22LSBOORCLXP1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSBOORCLXP1 0 0 ;
  SIZE 7.6 BY 3.6 ;
  SYMMETRY X Y ;
  SITE WCORE3600 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.117 LAYER MET1 ;
    ANTENNAMAXCUTCAR 25.643162 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 1 0.4 1.1 0.85 ;
        RECT 0.58 0.74 1.1 0.85 ;
      LAYER CUT01 ;
        RECT 0.625 0.745 0.715 0.835 ;
        RECT 1.005 0.45 1.095 0.54 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.0845 LAYER MET1 ;
    ANTENNAMAXCUTCAR 35.505803 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VYY ;
    PORT
      LAYER MET1 ;
        RECT 5.4 0.4 5.5 0.85 ;
        RECT 4.9 0.75 5.5 0.85 ;
      LAYER CUT01 ;
        RECT 4.945 0.755 5.035 0.845 ;
        RECT 5.405 0.45 5.495 0.54 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 1.245 2.82 ;
        RECT 7.1 0.78 8.1 2.82 ;
      LAYER MET1 ;
        RECT 0.075 1.595 0.255 1.96 ;
        RECT 0.095 1.64 0.275 2.005 ;
        RECT 0.395 1.64 0.575 2.005 ;
        RECT 0.635 1.595 0.815 1.96 ;
        RECT 0.955 1.64 1.135 2.005 ;
        RECT 0 1.64 7.6 1.96 ;
      LAYER CUT01 ;
        RECT 0.12 1.595 0.21 1.685 ;
        RECT 0.14 1.915 0.23 2.005 ;
        RECT 0.44 1.915 0.53 2.005 ;
        RECT 0.68 1.595 0.77 1.685 ;
        RECT 1 1.915 1.09 2.005 ;
        RECT 7.335 1.86 7.425 1.95 ;
        RECT 7.335 1.65 7.425 1.74 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.47 3.065 0.57 3.76 ;
        RECT 0.99 3.065 1.09 3.76 ;
        RECT 3.075 3.23 3.175 3.76 ;
        RECT 3.63 3.395 3.81 3.76 ;
        RECT 3.96 3.395 4.14 3.76 ;
        RECT 4.655 3.23 4.755 3.76 ;
        RECT 5.025 3.23 5.125 3.76 ;
        RECT 5.545 3.065 5.645 3.76 ;
        RECT 0 3.44 7.6 3.76 ;
        RECT 0.12 -0.16 0.22 0.535 ;
        RECT 0.64 -0.16 0.74 0.535 ;
        RECT 2.395 -0.16 2.495 0.56 ;
        RECT 2.93 -0.16 3.03 0.56 ;
        RECT 3.48 -0.16 3.58 0.56 ;
        RECT 4.015 -0.16 4.115 0.56 ;
        RECT 4.615 -0.16 4.715 0.43 ;
        RECT 5.135 -0.16 5.235 0.43 ;
        RECT 0 -0.16 7.6 0.16 ;
      LAYER CUT01 ;
        RECT 0.125 0.405 0.215 0.495 ;
        RECT 0.125 0.205 0.215 0.295 ;
        RECT 0.475 3.305 0.565 3.395 ;
        RECT 0.475 3.105 0.565 3.195 ;
        RECT 0.645 0.405 0.735 0.495 ;
        RECT 0.645 0.205 0.735 0.295 ;
        RECT 0.995 3.305 1.085 3.395 ;
        RECT 0.995 3.105 1.085 3.195 ;
        RECT 2.4 0.43 2.49 0.52 ;
        RECT 2.4 0.23 2.49 0.32 ;
        RECT 2.935 0.43 3.025 0.52 ;
        RECT 2.935 0.23 3.025 0.32 ;
        RECT 3.08 3.275 3.17 3.365 ;
        RECT 3.485 0.43 3.575 0.52 ;
        RECT 3.485 0.23 3.575 0.32 ;
        RECT 3.675 3.395 3.765 3.485 ;
        RECT 4.005 3.395 4.095 3.485 ;
        RECT 4.02 0.43 4.11 0.52 ;
        RECT 4.02 0.23 4.11 0.32 ;
        RECT 4.62 0.295 4.71 0.385 ;
        RECT 4.66 3.275 4.75 3.365 ;
        RECT 5.03 3.275 5.12 3.365 ;
        RECT 5.14 0.295 5.23 0.385 ;
        RECT 5.55 3.305 5.64 3.395 ;
        RECT 5.55 3.105 5.64 3.195 ;
    END
  END VSS
  PIN VYY
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT 2.245 0.78 6.1 2.82 ;
      LAYER MET1 ;
        RECT 0.06 2.125 7.54 2.275 ;
        RECT 2.395 1.14 2.495 1.475 ;
        RECT 4.555 1.14 4.655 1.475 ;
        RECT 5.85 1.14 5.95 1.475 ;
        RECT 0.06 1.325 7.54 1.475 ;
      LAYER CUT01 ;
        RECT 2.4 1.38 2.49 1.47 ;
        RECT 2.4 1.18 2.49 1.27 ;
        RECT 2.935 1.355 3.025 1.445 ;
        RECT 3.485 1.355 3.575 1.445 ;
        RECT 4.02 1.355 4.11 1.445 ;
        RECT 4.56 1.38 4.65 1.47 ;
        RECT 4.56 1.18 4.65 1.27 ;
        RECT 5.025 2.155 5.115 2.245 ;
        RECT 5.14 1.355 5.23 1.445 ;
        RECT 5.555 2.155 5.645 2.245 ;
        RECT 5.855 1.38 5.945 1.47 ;
        RECT 5.855 1.18 5.945 1.27 ;
    END
  END VYY
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.824 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 2.62 0.3 2.79 1.185 ;
        RECT 3.17 0.3 3.34 1.185 ;
        RECT 3.72 0.3 3.89 1.185 ;
        RECT 2.62 0.75 4.41 1.05 ;
        RECT 4.24 0.75 4.41 1.185 ;
      LAYER CUT01 ;
        RECT 2.66 1.075 2.75 1.165 ;
        RECT 2.66 0.505 2.75 0.595 ;
        RECT 2.66 0.305 2.75 0.395 ;
        RECT 3.21 1.075 3.3 1.165 ;
        RECT 3.21 0.505 3.3 0.595 ;
        RECT 3.21 0.305 3.3 0.395 ;
        RECT 3.76 1.075 3.85 1.165 ;
        RECT 3.76 0.505 3.85 0.595 ;
        RECT 3.76 0.305 3.85 0.395 ;
        RECT 4.28 1.075 4.37 1.165 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT 1.245 -0.5 2.245 4.1 ;
        RECT 6.1 -0.5 7.1 4.1 ;
        RECT -0.5 -0.5 8.1 0.78 ;
        RECT -0.5 2.82 8.1 4.1 ;
    END
  END VPW
  OBS
    LAYER MET1 ;
      RECT 0.38 0.285 0.48 1.225 ;
      RECT 1.26 0.4 1.36 1.225 ;
      RECT 0.335 1.125 1.36 1.225 ;
      RECT 0.685 2.375 0.875 2.475 ;
      RECT 0.73 2.8 1.415 2.9 ;
      RECT 2.87 2.975 4.355 3.075 ;
      RECT 1.315 2.8 1.415 3.28 ;
      RECT 2.87 2.975 2.97 3.28 ;
      RECT 1.315 3.18 2.97 3.28 ;
      RECT 0.73 2.375 0.83 3.315 ;
      RECT 1.985 2.375 2.565 2.475 ;
      RECT 2.665 2.775 4.8 2.875 ;
      RECT 1.985 2.375 2.085 3.08 ;
      RECT 2.665 2.775 2.765 3.08 ;
      RECT 1.985 2.98 2.765 3.08 ;
      RECT 2.185 2.575 5.385 2.675 ;
      RECT 4.455 3 5.385 3.1 ;
      RECT 4.455 3 4.555 3.275 ;
      RECT 3.335 3.175 4.555 3.275 ;
      RECT 5.285 2.575 5.385 3.315 ;
      RECT 4.875 0.4 4.975 0.64 ;
      RECT 4.7 0.54 4.975 0.64 ;
      RECT 4.7 0.54 4.8 1.05 ;
      RECT 4.7 0.95 4.975 1.05 ;
      RECT 4.875 0.95 4.975 1.225 ;
      RECT 4.875 1.125 5.485 1.225 ;
      RECT 2.87 2.375 5.955 2.475 ;
  END
END SC22LSBOORCLXP1

MACRO SC22LSDIANDCLXL1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSDIANDCLXL1 0 0 ;
  SIZE 3 BY 1.8 ;
  SYMMETRY X Y ;
  SITE CORE1800 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.181 LAYER MET1 ;
    ANTENNAMAXCUTCAR 42.556738 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.07 0.4 0.17 0.85 ;
        RECT 0.07 0.75 0.7 0.85 ;
        RECT 0.6 0.75 0.7 0.99 ;
        RECT 1.13 0.7 1.23 0.99 ;
        RECT 0.6 0.89 1.23 0.99 ;
      LAYER CUT01 ;
        RECT 0.075 0.45 0.165 0.54 ;
        RECT 0.435 0.75 0.525 0.84 ;
        RECT 1.135 0.74 1.225 0.83 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.1105 LAYER MET1 ;
    ANTENNAMAXCUTCAR 54.302862 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.31 0.4 0.41 0.65 ;
        RECT 0.31 0.55 0.92 0.65 ;
        RECT 0.82 0.5 0.92 0.79 ;
        RECT 0.82 0.5 1.43 0.6 ;
        RECT 1.33 0.5 1.43 0.79 ;
        RECT 1.33 0.69 1.67 0.79 ;
        RECT 1.57 0.69 1.67 0.875 ;
      LAYER CUT01 ;
        RECT 0.315 0.45 0.405 0.54 ;
        RECT 0.825 0.655 0.915 0.745 ;
        RECT 1.575 0.735 1.665 0.825 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.17 1.24 0.27 1.96 ;
        RECT 0.69 1.29 0.79 1.96 ;
        RECT 1.21 1.29 1.31 1.96 ;
        RECT 1.755 1.26 1.855 1.96 ;
        RECT 2.29 1.26 2.39 1.96 ;
        RECT 2.81 1.24 2.91 1.96 ;
        RECT 0 1.64 3 1.96 ;
      LAYER CUT01 ;
        RECT 0.175 1.5 0.265 1.59 ;
        RECT 0.175 1.28 0.265 1.37 ;
        RECT 0.695 1.53 0.785 1.62 ;
        RECT 0.695 1.33 0.785 1.42 ;
        RECT 1.215 1.53 1.305 1.62 ;
        RECT 1.215 1.33 1.305 1.42 ;
        RECT 1.76 1.5 1.85 1.59 ;
        RECT 1.76 1.3 1.85 1.39 ;
        RECT 2.295 1.5 2.385 1.59 ;
        RECT 2.295 1.3 2.385 1.39 ;
        RECT 2.815 1.5 2.905 1.59 ;
        RECT 2.815 1.28 2.905 1.37 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.71 -0.16 0.81 0.36 ;
        RECT 1.73 -0.16 1.83 0.36 ;
        RECT 2.25 -0.16 2.43 0.32 ;
        RECT 2.81 -0.16 2.91 0.555 ;
        RECT 0 -0.16 3 0.16 ;
      LAYER CUT01 ;
        RECT 0.715 0.225 0.805 0.315 ;
        RECT 1.735 0.225 1.825 0.315 ;
        RECT 2.295 0.225 2.385 0.315 ;
        RECT 2.815 0.425 2.905 0.515 ;
        RECT 2.815 0.225 2.905 0.315 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4372 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 1.995 0.96 2.165 1.295 ;
        RECT 1.995 0.44 2.685 0.6 ;
        RECT 2.485 0.44 2.685 1.12 ;
        RECT 1.995 0.96 2.685 1.12 ;
        RECT 2.515 0.44 2.685 1.295 ;
      LAYER CUT01 ;
        RECT 2.035 1.195 2.125 1.285 ;
        RECT 2.035 0.975 2.125 1.065 ;
        RECT 2.035 0.47 2.125 0.56 ;
        RECT 2.555 1.195 2.645 1.285 ;
        RECT 2.555 0.975 2.645 1.065 ;
        RECT 2.555 0.47 2.645 0.56 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT -0.5 -0.5 3.5 0.78 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 3.5 2.3 ;
    END
  END VNW
  OBS
    LAYER MET1 ;
      RECT 1.17 0.31 1.63 0.41 ;
      RECT 1.53 0.31 1.63 0.575 ;
      RECT 1.53 0.475 1.87 0.575 ;
      RECT 1.77 0.72 2.345 0.82 ;
      RECT 1.47 1 1.87 1.1 ;
      RECT 1.77 0.475 1.87 1.1 ;
      RECT 0.39 1.09 1.57 1.19 ;
      RECT 1.47 1 1.57 1.38 ;
      RECT 0.43 1.09 0.53 1.425 ;
      RECT 0.95 1.09 1.05 1.425 ;
  END
END SC22LSDIANDCLXL1

MACRO SC22LSDIANDCLXP1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSDIANDCLXP1 0 0 ;
  SIZE 4.8 BY 1.8 ;
  SYMMETRY X Y ;
  SITE CORE1800 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.28125 LAYER MET1 ;
    ANTENNAMAXCUTCAR 56.741946 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.07 0.4 0.17 0.85 ;
        RECT 0.07 0.75 0.8 0.85 ;
        RECT 0.7 0.75 0.8 1.05 ;
        RECT 1.35 0.7 1.45 1.05 ;
        RECT 2.31 0.69 2.41 1.05 ;
        RECT 0.7 0.95 2.41 1.05 ;
      LAYER CUT01 ;
        RECT 0.075 0.45 0.165 0.54 ;
        RECT 0.395 0.75 0.485 0.84 ;
        RECT 0.655 0.75 0.745 0.84 ;
        RECT 1.355 0.74 1.445 0.83 ;
        RECT 2.315 0.735 2.405 0.825 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.1755 LAYER MET1 ;
    ANTENNAMAXCUTCAR 51.286325 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.31 0.4 0.41 0.65 ;
        RECT 0.31 0.55 1.14 0.65 ;
        RECT 1.04 0.5 1.14 0.85 ;
        RECT 1.04 0.5 1.65 0.6 ;
        RECT 1.55 0.5 1.65 0.85 ;
        RECT 1.55 0.74 2.095 0.85 ;
      LAYER CUT01 ;
        RECT 0.315 0.45 0.405 0.54 ;
        RECT 1.045 0.72 1.135 0.81 ;
        RECT 1.955 0.74 2.045 0.83 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.39 1.4 0.49 1.96 ;
        RECT 0.91 1.4 1.01 1.96 ;
        RECT 1.43 1.4 1.53 1.96 ;
        RECT 1.95 1.4 2.05 1.96 ;
        RECT 2.5 1.4 2.6 1.96 ;
        RECT 3.05 1.25 3.15 1.96 ;
        RECT 3.57 1.24 3.67 1.96 ;
        RECT 4.09 1.24 4.19 1.96 ;
        RECT 4.61 1.24 4.71 1.96 ;
        RECT 0 1.64 4.8 1.96 ;
      LAYER CUT01 ;
        RECT 0.395 1.45 0.485 1.54 ;
        RECT 0.915 1.45 1.005 1.54 ;
        RECT 1.435 1.45 1.525 1.54 ;
        RECT 1.955 1.45 2.045 1.54 ;
        RECT 2.505 1.45 2.595 1.54 ;
        RECT 3.055 1.5 3.145 1.59 ;
        RECT 3.055 1.29 3.145 1.38 ;
        RECT 3.575 1.5 3.665 1.59 ;
        RECT 3.575 1.28 3.665 1.37 ;
        RECT 4.095 1.5 4.185 1.59 ;
        RECT 4.095 1.28 4.185 1.37 ;
        RECT 4.615 1.5 4.705 1.59 ;
        RECT 4.615 1.28 4.705 1.37 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.93 -0.16 1.03 0.36 ;
        RECT 1.95 -0.16 2.05 0.36 ;
        RECT 3.05 -0.16 3.15 0.57 ;
        RECT 3.57 -0.16 3.67 0.57 ;
        RECT 4.09 -0.16 4.19 0.57 ;
        RECT 4.61 -0.16 4.71 0.57 ;
        RECT 0 -0.16 4.8 0.16 ;
      LAYER CUT01 ;
        RECT 0.935 0.225 1.025 0.315 ;
        RECT 1.955 0.225 2.045 0.315 ;
        RECT 3.055 0.44 3.145 0.53 ;
        RECT 3.055 0.23 3.145 0.32 ;
        RECT 3.575 0.44 3.665 0.53 ;
        RECT 3.575 0.23 3.665 0.32 ;
        RECT 4.095 0.44 4.185 0.53 ;
        RECT 4.095 0.23 4.185 0.32 ;
        RECT 4.615 0.44 4.705 0.53 ;
        RECT 4.615 0.23 4.705 0.32 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.824 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 2.755 0.955 2.925 1.295 ;
        RECT 2.755 0.955 3.445 1.115 ;
        RECT 3.275 0.3 3.445 1.295 ;
        RECT 3.795 0.3 3.965 1.295 ;
        RECT 3.275 0.75 4.485 1.05 ;
        RECT 4.315 0.3 4.485 1.295 ;
      LAYER CUT01 ;
        RECT 2.795 1.195 2.885 1.285 ;
        RECT 2.795 0.975 2.885 1.065 ;
        RECT 3.315 1.195 3.405 1.285 ;
        RECT 3.315 0.975 3.405 1.065 ;
        RECT 3.315 0.505 3.405 0.595 ;
        RECT 3.315 0.305 3.405 0.395 ;
        RECT 3.835 1.195 3.925 1.285 ;
        RECT 3.835 0.975 3.925 1.065 ;
        RECT 3.835 0.505 3.925 0.595 ;
        RECT 3.835 0.305 3.925 0.395 ;
        RECT 4.355 1.195 4.445 1.285 ;
        RECT 4.355 0.975 4.445 1.065 ;
        RECT 4.355 0.505 4.445 0.595 ;
        RECT 4.355 0.305 4.445 0.395 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT -0.5 -0.5 5.3 0.78 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 5.3 2.3 ;
    END
  END VNW
  OBS
    LAYER MET1 ;
      RECT 1.39 0.31 1.85 0.41 ;
      RECT 1.75 0.31 1.85 0.575 ;
      RECT 1.75 0.475 2.615 0.575 ;
      RECT 2.515 0.715 3.135 0.815 ;
      RECT 2.515 0.475 2.615 1.25 ;
      RECT 0.13 1.15 2.615 1.25 ;
      RECT 0.13 1.01 0.23 1.385 ;
      RECT 0.65 1.15 0.75 1.485 ;
      RECT 1.17 1.15 1.27 1.485 ;
      RECT 1.69 1.15 1.79 1.485 ;
      RECT 2.21 1.15 2.31 1.485 ;
  END
END SC22LSDIANDCLXP1

MACRO SC22LSDICLXL1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSDICLXL1 0 0 ;
  SIZE 2.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE CORE1800 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.129 LAYER MET1 ;
    ANTENNAMAXCUTCAR 46.515202 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.07 0.4 0.17 0.85 ;
        RECT 0.07 0.74 0.815 0.85 ;
      LAYER CUT01 ;
        RECT 0.075 0.45 0.165 0.54 ;
        RECT 0.42 0.74 0.51 0.83 ;
        RECT 0.675 0.74 0.765 0.83 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.415 1.24 0.515 1.96 ;
        RECT 0.96 1.24 1.06 1.96 ;
        RECT 1.49 1.26 1.59 1.96 ;
        RECT 2.01 1.24 2.11 1.96 ;
        RECT 0 1.64 2.2 1.96 ;
      LAYER CUT01 ;
        RECT 0.42 1.5 0.51 1.59 ;
        RECT 0.42 1.28 0.51 1.37 ;
        RECT 0.965 1.5 1.055 1.59 ;
        RECT 0.965 1.28 1.055 1.37 ;
        RECT 1.495 1.5 1.585 1.59 ;
        RECT 1.495 1.3 1.585 1.39 ;
        RECT 2.015 1.5 2.105 1.59 ;
        RECT 2.015 1.28 2.105 1.37 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.675 -0.16 0.775 0.545 ;
        RECT 1.45 -0.16 1.63 0.32 ;
        RECT 2.01 -0.16 2.11 0.555 ;
        RECT 0 -0.16 2.2 0.16 ;
      LAYER CUT01 ;
        RECT 0.68 0.415 0.77 0.505 ;
        RECT 0.68 0.215 0.77 0.305 ;
        RECT 1.495 0.225 1.585 0.315 ;
        RECT 2.015 0.425 2.105 0.515 ;
        RECT 2.015 0.225 2.105 0.315 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4372 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 1.195 0.96 1.365 1.295 ;
        RECT 1.195 0.44 1.885 0.6 ;
        RECT 1.685 0.44 1.885 1.12 ;
        RECT 1.195 0.96 1.885 1.12 ;
        RECT 1.715 0.44 1.885 1.295 ;
      LAYER CUT01 ;
        RECT 1.235 1.195 1.325 1.285 ;
        RECT 1.235 0.975 1.325 1.065 ;
        RECT 1.235 0.47 1.325 0.56 ;
        RECT 1.755 1.195 1.845 1.285 ;
        RECT 1.755 0.975 1.845 1.065 ;
        RECT 1.755 0.47 1.845 0.56 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT -0.5 -0.5 2.7 0.78 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 2.7 2.3 ;
    END
  END VNW
  OBS
    LAYER MET1 ;
      RECT 0.935 0.72 1.545 0.82 ;
      RECT 0.935 0.285 1.035 1.09 ;
      RECT 0.155 0.99 1.035 1.09 ;
      RECT 0.675 0.99 0.775 1.335 ;
      RECT 0.155 0.99 0.255 1.375 ;
  END
END SC22LSDICLXL1

MACRO SC22LSDICLXP1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSDICLXP1 0 0 ;
  SIZE 4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE CORE1800 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.258 LAYER MET1 ;
    ANTENNAMAXCUTCAR 34.886494 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.07 0.4 0.17 0.85 ;
        RECT 0.07 0.73 1.01 0.85 ;
      LAYER CUT01 ;
        RECT 0.075 0.45 0.165 0.54 ;
        RECT 0.41 0.73 0.5 0.82 ;
        RECT 0.64 0.73 0.73 0.82 ;
        RECT 0.87 0.73 0.96 0.82 ;
    END
  END A
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.12 1.24 0.22 1.96 ;
        RECT 0.64 1.24 0.74 1.96 ;
        RECT 1.16 1.24 1.26 1.96 ;
        RECT 1.69 1.24 1.79 1.96 ;
        RECT 2.22 1.25 2.32 1.96 ;
        RECT 2.74 1.24 2.84 1.96 ;
        RECT 3.26 1.24 3.36 1.96 ;
        RECT 3.78 1.24 3.88 1.96 ;
        RECT 0 1.64 4 1.96 ;
      LAYER CUT01 ;
        RECT 0.125 1.5 0.215 1.59 ;
        RECT 0.125 1.28 0.215 1.37 ;
        RECT 0.645 1.5 0.735 1.59 ;
        RECT 0.645 1.28 0.735 1.37 ;
        RECT 1.165 1.5 1.255 1.59 ;
        RECT 1.165 1.28 1.255 1.37 ;
        RECT 1.695 1.5 1.785 1.59 ;
        RECT 1.695 1.28 1.785 1.37 ;
        RECT 2.225 1.5 2.315 1.59 ;
        RECT 2.225 1.29 2.315 1.38 ;
        RECT 2.745 1.5 2.835 1.59 ;
        RECT 2.745 1.28 2.835 1.37 ;
        RECT 3.265 1.5 3.355 1.59 ;
        RECT 3.265 1.28 3.355 1.37 ;
        RECT 3.785 1.5 3.875 1.59 ;
        RECT 3.785 1.28 3.875 1.37 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.9 -0.16 1 0.55 ;
        RECT 1.42 -0.16 1.52 0.55 ;
        RECT 2.22 -0.16 2.32 0.57 ;
        RECT 2.74 -0.16 2.84 0.57 ;
        RECT 3.26 -0.16 3.36 0.57 ;
        RECT 3.78 -0.16 3.88 0.57 ;
        RECT 0 -0.16 4 0.16 ;
      LAYER CUT01 ;
        RECT 0.905 0.42 0.995 0.51 ;
        RECT 0.905 0.21 0.995 0.3 ;
        RECT 1.425 0.42 1.515 0.51 ;
        RECT 1.425 0.21 1.515 0.3 ;
        RECT 2.225 0.44 2.315 0.53 ;
        RECT 2.225 0.23 2.315 0.32 ;
        RECT 2.745 0.44 2.835 0.53 ;
        RECT 2.745 0.23 2.835 0.32 ;
        RECT 3.265 0.44 3.355 0.53 ;
        RECT 3.265 0.23 3.355 0.32 ;
        RECT 3.785 0.44 3.875 0.53 ;
        RECT 3.785 0.23 3.875 0.32 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.824 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 1.925 0.955 2.095 1.295 ;
        RECT 1.925 0.955 2.615 1.115 ;
        RECT 2.445 0.3 2.615 1.295 ;
        RECT 2.965 0.3 3.135 1.295 ;
        RECT 2.445 0.75 3.655 1.05 ;
        RECT 3.485 0.3 3.655 1.295 ;
      LAYER CUT01 ;
        RECT 1.965 1.195 2.055 1.285 ;
        RECT 1.965 0.975 2.055 1.065 ;
        RECT 2.485 1.195 2.575 1.285 ;
        RECT 2.485 0.975 2.575 1.065 ;
        RECT 2.485 0.505 2.575 0.595 ;
        RECT 2.485 0.305 2.575 0.395 ;
        RECT 3.005 1.195 3.095 1.285 ;
        RECT 3.005 0.975 3.095 1.065 ;
        RECT 3.005 0.505 3.095 0.595 ;
        RECT 3.005 0.305 3.095 0.395 ;
        RECT 3.525 1.195 3.615 1.285 ;
        RECT 3.525 0.975 3.615 1.065 ;
        RECT 3.525 0.505 3.615 0.595 ;
        RECT 3.525 0.305 3.615 0.395 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT -0.5 -0.5 4.5 0.78 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 4.5 2.3 ;
    END
  END VNW
  OBS
    LAYER MET1 ;
      RECT 1.16 0.715 2.305 0.815 ;
      RECT 1.16 0.285 1.26 1.07 ;
      RECT 0.38 0.97 1.52 1.07 ;
      RECT 0.9 0.97 1 1.315 ;
      RECT 0.38 0.97 0.48 1.35 ;
      RECT 1.42 0.97 1.52 1.35 ;
  END
END SC22LSDICLXP1

MACRO SC22LSDIORCLXL1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSDIORCLXL1 0 0 ;
  SIZE 4.2 BY 1.8 ;
  SYMMETRY X Y ;
  SITE CORE1800 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.20425 LAYER MET1 ;
    ANTENNAMAXCUTCAR 47.434535 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.825 0.4 0.925 0.85 ;
        RECT 1.745 0.55 1.845 0.85 ;
        RECT 0.825 0.55 2.6 0.65 ;
        RECT 2.5 0.55 2.6 0.8 ;
        RECT 2.5 0.7 2.865 0.8 ;
      LAYER CUT01 ;
        RECT 0.83 0.72 0.92 0.81 ;
        RECT 0.83 0.455 0.92 0.545 ;
        RECT 1.75 0.715 1.84 0.805 ;
        RECT 2.73 0.705 2.82 0.795 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.05725 LAYER MET1 ;
    ANTENNAMAXCUTCAR 52.406044 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.1 0.325 0.2 0.85 ;
        RECT 0.1 0.75 0.305 0.85 ;
        RECT 0.1 0.325 0.725 0.415 ;
      LAYER CUT01 ;
        RECT 0.165 0.755 0.255 0.845 ;
        RECT 0.585 0.325 0.675 0.415 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.345 1.25 0.445 1.96 ;
        RECT 1.28 1.4 1.38 1.96 ;
        RECT 2.21 1.4 2.31 1.96 ;
        RECT 2.98 1.25 3.08 1.96 ;
        RECT 3.5 1.26 3.6 1.96 ;
        RECT 4.02 1.24 4.12 1.96 ;
        RECT 0 1.64 4.2 1.96 ;
      LAYER CUT01 ;
        RECT 0.35 1.5 0.44 1.59 ;
        RECT 0.35 1.29 0.44 1.38 ;
        RECT 1.285 1.45 1.375 1.54 ;
        RECT 2.215 1.45 2.305 1.54 ;
        RECT 2.985 1.5 3.075 1.59 ;
        RECT 2.985 1.29 3.075 1.38 ;
        RECT 3.505 1.5 3.595 1.59 ;
        RECT 3.505 1.3 3.595 1.39 ;
        RECT 4.025 1.5 4.115 1.59 ;
        RECT 4.025 1.28 4.115 1.37 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.075 -0.16 0.175 0.225 ;
        RECT 1.95 -0.16 2.05 0.38 ;
        RECT 2.435 -0.16 2.615 0.23 ;
        RECT 3 -0.16 3.1 0.38 ;
        RECT 3.46 -0.16 3.64 0.32 ;
        RECT 4.02 -0.16 4.12 0.555 ;
        RECT 0 -0.16 4.2 0.16 ;
      LAYER CUT01 ;
        RECT 0.08 0.095 0.17 0.185 ;
        RECT 1.955 0.245 2.045 0.335 ;
        RECT 2.48 0.14 2.57 0.23 ;
        RECT 3.005 0.245 3.095 0.335 ;
        RECT 3.505 0.225 3.595 0.315 ;
        RECT 4.025 0.425 4.115 0.515 ;
        RECT 4.025 0.225 4.115 0.315 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.4372 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 3.205 0.96 3.375 1.295 ;
        RECT 3.205 0.44 3.895 0.6 ;
        RECT 3.695 0.44 3.895 1.12 ;
        RECT 3.205 0.96 3.895 1.12 ;
        RECT 3.725 0.44 3.895 1.295 ;
      LAYER CUT01 ;
        RECT 3.245 1.195 3.335 1.285 ;
        RECT 3.245 0.975 3.335 1.065 ;
        RECT 3.245 0.47 3.335 0.56 ;
        RECT 3.765 1.195 3.855 1.285 ;
        RECT 3.765 0.975 3.855 1.065 ;
        RECT 3.765 0.47 3.855 0.56 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT -0.5 -0.5 4.7 0.78 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 4.7 2.3 ;
    END
  END VNW
  OBS
    LAYER MET1 ;
      RECT 0.3 0.505 0.55 0.605 ;
      RECT 1.235 0.75 1.425 0.85 ;
      RECT 2.1 0.75 2.355 0.85 ;
      RECT 0.45 0.505 0.55 1.05 ;
      RECT 1.28 0.75 1.38 1.05 ;
      RECT 2.1 0.75 2.2 1.05 ;
      RECT 0.08 0.95 2.2 1.05 ;
      RECT 0.08 0.95 0.18 1.325 ;
      RECT 2.17 0.35 2.88 0.45 ;
      RECT 2.78 0.35 2.88 0.59 ;
      RECT 2.78 0.49 3.075 0.59 ;
      RECT 2.975 0.72 3.555 0.82 ;
      RECT 2.975 0.49 3.075 1.05 ;
      RECT 2.74 0.95 3.075 1.05 ;
      RECT 0.775 1.15 2.84 1.25 ;
      RECT 2.74 0.95 2.84 1.39 ;
      RECT 0.815 1.15 0.915 1.485 ;
      RECT 1.745 1.15 1.845 1.485 ;
  END
END SC22LSDIORCLXL1

MACRO SC22LSDIORCLXP1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN SC22LSDIORCLXP1 0 0 ;
  SIZE 6.4 BY 1.8 ;
  SYMMETRY X Y ;
  SITE CORE1800 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.29325 LAYER MET1 ;
    ANTENNAMAXCUTCAR 59.118062 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 1.11 0.4 1.21 0.85 ;
        RECT 2.01 0.55 2.11 0.85 ;
        RECT 3 0.55 3.1 0.83 ;
        RECT 1.11 0.55 3.72 0.65 ;
        RECT 3.62 0.55 3.72 0.785 ;
        RECT 3.62 0.685 3.92 0.785 ;
        RECT 3.82 0.685 3.92 0.875 ;
      LAYER CUT01 ;
        RECT 1.115 0.72 1.205 0.81 ;
        RECT 1.115 0.445 1.205 0.535 ;
        RECT 2.015 0.715 2.105 0.805 ;
        RECT 3.005 0.69 3.095 0.78 ;
        RECT 3.825 0.735 3.915 0.825 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNAGATEAREA 0.117 LAYER MET1 ;
    ANTENNAMAXCUTCAR 25.643162 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDD ;
    PORT
      LAYER MET1 ;
        RECT 0.53 0.35 0.63 0.85 ;
        RECT 0.3 0.74 0.63 0.85 ;
        RECT 0.53 0.35 1.01 0.45 ;
      LAYER CUT01 ;
        RECT 0.35 0.74 0.44 0.83 ;
        RECT 0.875 0.355 0.965 0.445 ;
    END
  END EN
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.07 1.25 0.17 1.96 ;
        RECT 0.61 1.25 0.71 1.96 ;
        RECT 1.55 1.4 1.65 1.96 ;
        RECT 2.47 1.4 2.57 1.96 ;
        RECT 3.46 1.4 3.56 1.96 ;
        RECT 4.15 1.25 4.25 1.96 ;
        RECT 4.67 1.25 4.77 1.96 ;
        RECT 5.19 1.24 5.29 1.96 ;
        RECT 5.71 1.24 5.81 1.96 ;
        RECT 6.23 1.24 6.33 1.96 ;
        RECT 0 1.64 6.4 1.96 ;
      LAYER CUT01 ;
        RECT 0.075 1.5 0.165 1.59 ;
        RECT 0.075 1.29 0.165 1.38 ;
        RECT 0.615 1.5 0.705 1.59 ;
        RECT 0.615 1.29 0.705 1.38 ;
        RECT 1.555 1.45 1.645 1.54 ;
        RECT 2.475 1.45 2.565 1.54 ;
        RECT 3.465 1.45 3.555 1.54 ;
        RECT 4.155 1.5 4.245 1.59 ;
        RECT 4.155 1.29 4.245 1.38 ;
        RECT 4.675 1.5 4.765 1.59 ;
        RECT 4.675 1.29 4.765 1.38 ;
        RECT 5.195 1.5 5.285 1.59 ;
        RECT 5.195 1.28 5.285 1.37 ;
        RECT 5.715 1.5 5.805 1.59 ;
        RECT 5.715 1.28 5.805 1.37 ;
        RECT 6.235 1.5 6.325 1.59 ;
        RECT 6.235 1.28 6.325 1.37 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.07 -0.16 0.17 0.365 ;
        RECT 0.625 -0.16 0.725 0.25 ;
        RECT 2.21 -0.16 2.31 0.375 ;
        RECT 2.695 -0.16 2.875 0.23 ;
        RECT 3.32 -0.16 3.5 0.23 ;
        RECT 4.02 -0.16 4.12 0.375 ;
        RECT 4.67 -0.16 4.77 0.57 ;
        RECT 5.19 -0.16 5.29 0.57 ;
        RECT 5.71 -0.16 5.81 0.57 ;
        RECT 6.23 -0.16 6.33 0.57 ;
        RECT 0 -0.16 6.4 0.16 ;
      LAYER CUT01 ;
        RECT 0.075 0.225 0.165 0.315 ;
        RECT 0.63 0.115 0.72 0.205 ;
        RECT 2.215 0.24 2.305 0.33 ;
        RECT 2.74 0.14 2.83 0.23 ;
        RECT 3.365 0.14 3.455 0.23 ;
        RECT 4.025 0.24 4.115 0.33 ;
        RECT 4.675 0.44 4.765 0.53 ;
        RECT 4.675 0.23 4.765 0.32 ;
        RECT 5.195 0.44 5.285 0.53 ;
        RECT 5.195 0.23 5.285 0.32 ;
        RECT 5.715 0.44 5.805 0.53 ;
        RECT 5.715 0.23 5.805 0.32 ;
        RECT 6.235 0.44 6.325 0.53 ;
        RECT 6.235 0.23 6.325 0.32 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.824 LAYER MET1 ;
    PORT
      LAYER MET1 ;
        RECT 4.375 0.955 4.545 1.295 ;
        RECT 4.375 0.955 5.065 1.115 ;
        RECT 4.895 0.3 5.065 1.295 ;
        RECT 5.415 0.3 5.585 1.295 ;
        RECT 4.895 0.75 6.105 1.05 ;
        RECT 5.935 0.3 6.105 1.295 ;
      LAYER CUT01 ;
        RECT 4.415 1.195 4.505 1.285 ;
        RECT 4.415 0.975 4.505 1.065 ;
        RECT 4.935 1.195 5.025 1.285 ;
        RECT 4.935 0.975 5.025 1.065 ;
        RECT 4.935 0.505 5.025 0.595 ;
        RECT 4.935 0.305 5.025 0.395 ;
        RECT 5.455 1.195 5.545 1.285 ;
        RECT 5.455 0.975 5.545 1.065 ;
        RECT 5.455 0.505 5.545 0.595 ;
        RECT 5.455 0.305 5.545 0.395 ;
        RECT 5.975 1.195 6.065 1.285 ;
        RECT 5.975 0.975 6.065 1.065 ;
        RECT 5.975 0.505 6.065 0.595 ;
        RECT 5.975 0.305 6.065 0.395 ;
    END
  END Y
  PIN VPW
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER PWELL ;
        RECT -0.5 -0.5 6.9 0.78 ;
    END
  END VPW
  PIN VNW
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER NWELL ;
        RECT -0.5 0.78 6.9 2.3 ;
    END
  END VNW
  OBS
    LAYER MET1 ;
      RECT 0.33 0.41 0.43 0.61 ;
      RECT 0.1 0.51 0.43 0.61 ;
      RECT 1.505 0.75 1.695 0.85 ;
      RECT 2.425 0.75 2.615 0.85 ;
      RECT 3.285 0.75 3.52 0.85 ;
      RECT 0.1 0.51 0.2 1.05 ;
      RECT 0.73 0.675 0.83 1.05 ;
      RECT 1.55 0.75 1.65 1.05 ;
      RECT 2.47 0.75 2.57 1.05 ;
      RECT 3.285 0.75 3.385 1.05 ;
      RECT 0.1 0.95 3.385 1.05 ;
      RECT 0.33 0.95 0.43 1.32 ;
      RECT 2.43 0.35 3.92 0.45 ;
      RECT 3.82 0.35 3.92 0.585 ;
      RECT 3.82 0.485 4.14 0.585 ;
      RECT 4.04 0.715 4.755 0.815 ;
      RECT 4.04 0.485 4.14 1.11 ;
      RECT 3.92 1.01 4.14 1.11 ;
      RECT 1.05 1.15 4.02 1.25 ;
      RECT 3.92 1.01 4.02 1.44 ;
      RECT 1.09 1.15 1.19 1.485 ;
      RECT 2.01 1.15 2.11 1.485 ;
      RECT 3 1.15 3.1 1.485 ;
  END
END SC22LSDIORCLXP1

END LIBRARY
VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
#
#   MOL INFORMATION (TECH)
#       SCHEMA : 02/05/08 (V=107)
#       CARD   : 06/02/03 (V=1)
#
#
#   MOL INFORMATION (PC)
#       SCHEMA : 02/05/08 (V=107)
#       CARD   : 07/07/27 (V=1)
#
#MACRO SECTION
  MACRO RAM200
    CLASS BLOCK ;
    FOREIGN RAM200  0.000 0.000 ;
    SIZE 84.395 BY 188.535 ;
    SYMMETRY R90 X Y ;
    PIN IA[9]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 12.175 0.000 12.275 0.380 ;
          LAYER MET2 ;
          RECT 12.175 0.000 12.275 0.380 ;
      END
    END IA[9]
    PIN IA[8]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 27.230 0.000 27.330 0.380 ;
          LAYER MET2 ;
          RECT 27.230 0.000 27.330 0.380 ;
      END
    END IA[8]
    PIN IA[7]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 25.785 0.000 25.885 0.380 ;
          LAYER MET2 ;
          RECT 25.785 0.000 25.885 0.380 ;
      END
    END IA[7]
    PIN IA[6]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 24.340 0.000 24.440 0.380 ;
          LAYER MET2 ;
          RECT 24.340 0.000 24.440 0.380 ;
      END
    END IA[6]
    PIN IA[5]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 22.895 0.000 22.995 0.380 ;
          LAYER MET2 ;
          RECT 22.895 0.000 22.995 0.380 ;
      END
    END IA[5]
    PIN IA[4]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 21.450 0.000 21.550 0.380 ;
          LAYER MET2 ;
          RECT 21.450 0.000 21.550 0.380 ;
      END
    END IA[4]
    PIN IA[3]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 20.005 0.000 20.105 0.380 ;
          LAYER MET2 ;
          RECT 20.005 0.000 20.105 0.380 ;
      END
    END IA[3]
    PIN IA[2]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 17.955 0.000 18.055 0.380 ;
          LAYER MET2 ;
          RECT 17.955 0.000 18.055 0.380 ;
      END
    END IA[2]
    PIN IA[1]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 16.510 0.000 16.610 0.380 ;
          LAYER MET2 ;
          RECT 16.510 0.000 16.610 0.380 ;
      END
    END IA[1]
    PIN IA[0]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 15.065 0.000 15.165 0.380 ;
          LAYER MET2 ;
          RECT 15.065 0.000 15.165 0.380 ;
      END
    END IA[0]
    PIN BP
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 2.490 0.000 2.590 0.380 ;
          LAYER MET2 ;
          RECT 2.490 0.000 2.590 0.380 ;
      END
    END BP
    PIN WE
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 30.120 0.000 30.220 0.380 ;
          LAYER MET2 ;
          RECT 30.120 0.000 30.220 0.380 ;
      END
    END WE
    PIN CE
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 6.680 0.000 6.780 0.380 ;
          LAYER MET2 ;
          RECT 6.680 0.000 6.780 0.380 ;
      END
    END CE
    PIN CK
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 5.800 0.000 5.900 0.380 ;
          LAYER MET2 ;
          RECT 5.800 0.000 5.900 0.380 ;
      END
    END CK
    PIN A[9]
      DIRECTION OUTPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 81.315 0.000 81.415 0.380 ;
          LAYER MET2 ;
          RECT 81.315 0.000 81.415 0.380 ;
      END
    END A[9]
    PIN I[9]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 78.715 0.000 78.815 0.380 ;
          LAYER MET2 ;
          RECT 78.715 0.000 78.815 0.380 ;
      END
    END I[9]
    PIN DM[9]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 79.475 0.000 79.575 0.380 ;
          LAYER MET2 ;
          RECT 79.475 0.000 79.575 0.380 ;
      END
    END DM[9]
    PIN A[8]
      DIRECTION OUTPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 77.195 0.000 77.295 0.380 ;
          LAYER MET2 ;
          RECT 77.195 0.000 77.295 0.380 ;
      END
    END A[8]
    PIN I[8]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 74.595 0.000 74.695 0.380 ;
          LAYER MET2 ;
          RECT 74.595 0.000 74.695 0.380 ;
      END
    END I[8]
    PIN DM[8]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 75.355 0.000 75.455 0.380 ;
          LAYER MET2 ;
          RECT 75.355 0.000 75.455 0.380 ;
      END
    END DM[8]
    PIN A[7]
      DIRECTION OUTPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 73.075 0.000 73.175 0.380 ;
          LAYER MET2 ;
          RECT 73.075 0.000 73.175 0.380 ;
      END
    END A[7]
    PIN I[7]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 70.475 0.000 70.575 0.380 ;
          LAYER MET2 ;
          RECT 70.475 0.000 70.575 0.380 ;
      END
    END I[7]
    PIN DM[7]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 71.235 0.000 71.335 0.380 ;
          LAYER MET2 ;
          RECT 71.235 0.000 71.335 0.380 ;
      END
    END DM[7]
    PIN A[6]
      DIRECTION OUTPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 68.955 0.000 69.055 0.380 ;
          LAYER MET2 ;
          RECT 68.955 0.000 69.055 0.380 ;
      END
    END A[6]
    PIN I[6]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 66.355 0.000 66.455 0.380 ;
          LAYER MET2 ;
          RECT 66.355 0.000 66.455 0.380 ;
      END
    END I[6]
    PIN DM[6]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 67.115 0.000 67.215 0.380 ;
          LAYER MET2 ;
          RECT 67.115 0.000 67.215 0.380 ;
      END
    END DM[6]
    PIN A[5]
      DIRECTION OUTPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 64.835 0.000 64.935 0.380 ;
          LAYER MET2 ;
          RECT 64.835 0.000 64.935 0.380 ;
      END
    END A[5]
    PIN I[5]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 62.235 0.000 62.335 0.380 ;
          LAYER MET2 ;
          RECT 62.235 0.000 62.335 0.380 ;
      END
    END I[5]
    PIN DM[5]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 62.995 0.000 63.095 0.380 ;
          LAYER MET2 ;
          RECT 62.995 0.000 63.095 0.380 ;
      END
    END DM[5]
    PIN A[4]
      DIRECTION OUTPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 60.715 0.000 60.815 0.380 ;
          LAYER MET2 ;
          RECT 60.715 0.000 60.815 0.380 ;
      END
    END A[4]
    PIN I[4]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 58.115 0.000 58.215 0.380 ;
          LAYER MET2 ;
          RECT 58.115 0.000 58.215 0.380 ;
      END
    END I[4]
    PIN DM[4]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 58.875 0.000 58.975 0.380 ;
          LAYER MET2 ;
          RECT 58.875 0.000 58.975 0.380 ;
      END
    END DM[4]
    PIN A[3]
      DIRECTION OUTPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 56.595 0.000 56.695 0.380 ;
          LAYER MET2 ;
          RECT 56.595 0.000 56.695 0.380 ;
      END
    END A[3]
    PIN I[3]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 53.995 0.000 54.095 0.380 ;
          LAYER MET2 ;
          RECT 53.995 0.000 54.095 0.380 ;
      END
    END I[3]
    PIN DM[3]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 54.755 0.000 54.855 0.380 ;
          LAYER MET2 ;
          RECT 54.755 0.000 54.855 0.380 ;
      END
    END DM[3]
    PIN A[2]
      DIRECTION OUTPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 52.475 0.000 52.575 0.380 ;
          LAYER MET2 ;
          RECT 52.475 0.000 52.575 0.380 ;
      END
    END A[2]
    PIN I[2]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 49.875 0.000 49.975 0.380 ;
          LAYER MET2 ;
          RECT 49.875 0.000 49.975 0.380 ;
      END
    END I[2]
    PIN DM[2]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 50.635 0.000 50.735 0.380 ;
          LAYER MET2 ;
          RECT 50.635 0.000 50.735 0.380 ;
      END
    END DM[2]
    PIN A[1]
      DIRECTION OUTPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 48.355 0.000 48.455 0.380 ;
          LAYER MET2 ;
          RECT 48.355 0.000 48.455 0.380 ;
      END
    END A[1]
    PIN I[1]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 45.755 0.000 45.855 0.380 ;
          LAYER MET2 ;
          RECT 45.755 0.000 45.855 0.380 ;
      END
    END I[1]
    PIN DM[1]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 46.515 0.000 46.615 0.380 ;
          LAYER MET2 ;
          RECT 46.515 0.000 46.615 0.380 ;
      END
    END DM[1]
    PIN A[0]
      DIRECTION OUTPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 44.235 0.000 44.335 0.380 ;
          LAYER MET2 ;
          RECT 44.235 0.000 44.335 0.380 ;
      END
    END A[0]
    PIN I[0]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 41.635 0.000 41.735 0.380 ;
          LAYER MET2 ;
          RECT 41.635 0.000 41.735 0.380 ;
      END
    END I[0]
    PIN DM[0]
      DIRECTION INPUT ;
      USE SIGNAL ;
      ANTENNADIFFAREA 0.100 ;
      PORT
          LAYER MET3 ;
          RECT 42.395 0.000 42.495 0.380 ;
          LAYER MET2 ;
          RECT 42.395 0.000 42.495 0.380 ;
      END
    END DM[0]
    PIN VDD
      DIRECTION INOUT ;
      USE POWER ;
      SHAPE ABUTMENT ;
      PORT
          LAYER MET4 ;
          RECT 43.330 1.500 43.930 185.970 ;
          LAYER MET4 ;
          RECT 47.450 1.500 48.050 185.970 ;
          LAYER MET4 ;
          RECT 51.570 1.500 52.170 185.970 ;
          LAYER MET4 ;
          RECT 55.690 1.500 56.290 185.970 ;
          LAYER MET4 ;
          RECT 59.810 1.500 60.410 185.970 ;
          LAYER MET4 ;
          RECT 63.930 1.500 64.530 185.970 ;
          LAYER MET4 ;
          RECT 68.050 1.500 68.650 185.970 ;
          LAYER MET4 ;
          RECT 72.170 1.500 72.770 185.970 ;
          LAYER MET4 ;
          RECT 76.290 1.500 76.890 185.970 ;
          LAYER MET4 ;
          RECT 80.410 1.500 81.010 185.970 ;
          LAYER MET4 ;
          RECT 3.050 1.500 4.550 186.050 ;
          LAYER MET4 ;
          RECT 9.290 1.500 10.790 186.050 ;
          LAYER MET4 ;
          RECT 15.530 1.500 17.030 186.050 ;
          LAYER MET4 ;
          RECT 22.380 1.500 23.880 186.050 ;
          LAYER MET4 ;
          RECT 28.620 1.500 30.120 186.050 ;
          LAYER MET4 ;
          RECT 34.860 1.500 36.360 186.050 ;
      END
    END VDD
    PIN VSS
      DIRECTION INOUT ;
      USE GROUND ;
      SHAPE ABUTMENT ;
      PORT
          LAYER MET4 ;
          RECT 41.270 1.500 41.870 185.970 ;
          LAYER MET4 ;
          RECT 45.390 1.500 45.990 185.970 ;
          LAYER MET4 ;
          RECT 49.510 1.500 50.110 185.970 ;
          LAYER MET4 ;
          RECT 53.630 1.500 54.230 185.970 ;
          LAYER MET4 ;
          RECT 57.750 1.500 58.350 185.970 ;
          LAYER MET4 ;
          RECT 61.870 1.500 62.470 185.970 ;
          LAYER MET4 ;
          RECT 65.990 1.500 66.590 185.970 ;
          LAYER MET4 ;
          RECT 70.110 1.500 70.710 185.970 ;
          LAYER MET4 ;
          RECT 74.230 1.500 74.830 185.970 ;
          LAYER MET4 ;
          RECT 78.350 1.500 78.950 185.970 ;
          LAYER MET4 ;
          RECT 6.170 1.500 7.670 186.050 ;
          LAYER MET4 ;
          RECT 12.410 1.500 13.910 186.050 ;
          LAYER MET4 ;
          RECT 19.260 1.500 20.760 186.050 ;
          LAYER MET4 ;
          RECT 25.500 1.500 27.000 186.050 ;
          LAYER MET4 ;
          RECT 31.740 1.500 33.240 186.050 ;
      END
    END VSS
    OBS
      LAYER MET1 ;
      RECT 0.000 0.000 84.395 188.535 ;
      LAYER CUT12 ;
      RECT 0.000 0.000 84.395 188.535 ;
      LAYER MET2 ;
      RECT 0.000 0.000 84.395 188.535 ;
      LAYER CUT23 ;
      RECT 0.000 0.000 84.395 188.535 ;
      LAYER MET3 ;
      RECT 0.000 0.000 84.395 188.535 ;
      LAYER CUT34 ;
      RECT 0.000 0.000 84.395 188.535 ;
      LAYER MET4 ;
      RECT 0.000 0.000 84.395 188.535 ;
    END
  END RAM200
END LIBRARY
#------------------------------------------------------------------
# cs202_pgpsw.lef
# designed by FVD)DSIpj
#
# Rev. 3.0  2007/09/13  added DSIPGX2LBFC1, DSIPGX2LBFF1, DSIPGX2LBFJ1,
#                       DSIPGX2LBFL1, DSIPGX2LBFN1, DSIPGX2LCNRC2,
#                       DSIPGX2LPSRCS2, DSIPGX2LSPRCS2
#                       defined "SHAPE ABUTMENT" in each power pin
#                       GDS: cs202_pgpsw.gds(Rev. 3.0)
# Rev. 2.0  2007/07/04  added DSIPGX2LCNRC1
#                       GDS: cs202_pgpsw.gds(Rev. 2.0)
# Rev. 1.0  2007/06/15  new release
#                       GDS: cs202_pgpsw.gds(Rev. 1.0)
#------------------------------------------------------------------

VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

SITE CORE1800
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 0.200 BY 1.800 ;
END CORE1800

SITE WCORE3600
  CLASS CORE ;
  SYMMETRY X Y ;
  SIZE 0.200 BY 3.600 ;
END WCORE3600

MACRO DSIPGX2LBFC1
  CLASS RING ;
  ORIGIN 0 0 ;
  FOREIGN DSIPGX2LBFC1 0 0 ;
  SIZE 11.57 BY 11.57 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.23 0.23 0.37 11.57 ;
        RECT 0.23 0.23 11.57 0.37 ;
      LAYER CUT01 ;
        RECT 0.255 11.255 0.345 11.345 ;
        RECT 0.255 11.035 0.345 11.125 ;
        RECT 0.255 10.815 0.345 10.905 ;
        RECT 0.255 10.595 0.345 10.685 ;
        RECT 0.255 10.375 0.345 10.465 ;
        RECT 0.255 10.155 0.345 10.245 ;
        RECT 0.255 9.935 0.345 10.025 ;
        RECT 0.255 9.715 0.345 9.805 ;
        RECT 0.255 9.495 0.345 9.585 ;
        RECT 0.255 9.275 0.345 9.365 ;
        RECT 0.255 9.055 0.345 9.145 ;
        RECT 0.255 8.835 0.345 8.925 ;
        RECT 0.255 8.615 0.345 8.705 ;
        RECT 0.255 8.395 0.345 8.485 ;
        RECT 0.255 8.175 0.345 8.265 ;
        RECT 0.255 7.955 0.345 8.045 ;
        RECT 0.255 7.735 0.345 7.825 ;
        RECT 0.255 7.515 0.345 7.605 ;
        RECT 0.255 7.295 0.345 7.385 ;
        RECT 0.255 7.075 0.345 7.165 ;
        RECT 0.255 6.855 0.345 6.945 ;
        RECT 0.255 6.635 0.345 6.725 ;
        RECT 0.255 6.415 0.345 6.505 ;
        RECT 0.255 6.195 0.345 6.285 ;
        RECT 0.255 5.975 0.345 6.065 ;
        RECT 0.255 5.755 0.345 5.845 ;
        RECT 0.255 5.535 0.345 5.625 ;
        RECT 0.255 5.315 0.345 5.405 ;
        RECT 0.255 5.095 0.345 5.185 ;
        RECT 0.255 4.875 0.345 4.965 ;
        RECT 0.255 4.655 0.345 4.745 ;
        RECT 0.255 4.435 0.345 4.525 ;
        RECT 0.255 4.215 0.345 4.305 ;
        RECT 0.255 3.995 0.345 4.085 ;
        RECT 0.255 3.775 0.345 3.865 ;
        RECT 0.255 3.555 0.345 3.645 ;
        RECT 0.255 3.335 0.345 3.425 ;
        RECT 0.255 3.115 0.345 3.205 ;
        RECT 0.255 2.895 0.345 2.985 ;
        RECT 0.255 2.675 0.345 2.765 ;
        RECT 0.255 2.455 0.345 2.545 ;
        RECT 0.255 2.235 0.345 2.325 ;
        RECT 0.255 2.015 0.345 2.105 ;
        RECT 0.255 1.795 0.345 1.885 ;
        RECT 0.255 1.575 0.345 1.665 ;
        RECT 0.255 1.355 0.345 1.445 ;
        RECT 0.255 1.135 0.345 1.225 ;
        RECT 0.255 0.915 0.345 1.005 ;
        RECT 0.255 0.695 0.345 0.785 ;
        RECT 0.255 0.475 0.345 0.565 ;
        RECT 0.475 0.255 0.565 0.345 ;
        RECT 0.695 0.255 0.785 0.345 ;
        RECT 0.915 0.255 1.005 0.345 ;
        RECT 1.135 0.255 1.225 0.345 ;
        RECT 1.355 0.255 1.445 0.345 ;
        RECT 1.575 0.255 1.665 0.345 ;
        RECT 1.795 0.255 1.885 0.345 ;
        RECT 2.015 0.255 2.105 0.345 ;
        RECT 2.235 0.255 2.325 0.345 ;
        RECT 2.455 0.255 2.545 0.345 ;
        RECT 2.675 0.255 2.765 0.345 ;
        RECT 2.895 0.255 2.985 0.345 ;
        RECT 3.115 0.255 3.205 0.345 ;
        RECT 3.335 0.255 3.425 0.345 ;
        RECT 3.555 0.255 3.645 0.345 ;
        RECT 3.775 0.255 3.865 0.345 ;
        RECT 3.995 0.255 4.085 0.345 ;
        RECT 4.215 0.255 4.305 0.345 ;
        RECT 4.435 0.255 4.525 0.345 ;
        RECT 4.655 0.255 4.745 0.345 ;
        RECT 4.875 0.255 4.965 0.345 ;
        RECT 5.095 0.255 5.185 0.345 ;
        RECT 5.315 0.255 5.405 0.345 ;
        RECT 5.535 0.255 5.625 0.345 ;
        RECT 5.755 0.255 5.845 0.345 ;
        RECT 5.975 0.255 6.065 0.345 ;
        RECT 6.195 0.255 6.285 0.345 ;
        RECT 6.415 0.255 6.505 0.345 ;
        RECT 6.635 0.255 6.725 0.345 ;
        RECT 6.855 0.255 6.945 0.345 ;
        RECT 7.075 0.255 7.165 0.345 ;
        RECT 7.295 0.255 7.385 0.345 ;
        RECT 7.515 0.255 7.605 0.345 ;
        RECT 7.735 0.255 7.825 0.345 ;
        RECT 7.955 0.255 8.045 0.345 ;
        RECT 8.175 0.255 8.265 0.345 ;
        RECT 8.395 0.255 8.485 0.345 ;
        RECT 8.615 0.255 8.705 0.345 ;
        RECT 8.835 0.255 8.925 0.345 ;
        RECT 9.055 0.255 9.145 0.345 ;
        RECT 9.275 0.255 9.365 0.345 ;
        RECT 9.495 0.255 9.585 0.345 ;
        RECT 9.715 0.255 9.805 0.345 ;
        RECT 9.935 0.255 10.025 0.345 ;
        RECT 10.155 0.255 10.245 0.345 ;
        RECT 10.375 0.255 10.465 0.345 ;
        RECT 10.595 0.255 10.685 0.345 ;
        RECT 10.815 0.255 10.905 0.345 ;
        RECT 11.035 0.255 11.125 0.345 ;
        RECT 11.255 0.255 11.345 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 0.036 LAYER MET1 ;
      ANTENNAGATEAREA 0.036 LAYER MET2 ;
    ANTENNAMAXCUTCAR 416.666667 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDDSRC ;
    PORT
      LAYER CUT01 ;
        RECT 2.345 5.905 2.435 5.995 ;
      LAYER MET1 ;
        RECT 1.855 5.415 1.955 6 ;
        RECT 1.855 5.9 2.44 6 ;
        RECT 2.34 5.865 2.44 6.035 ;
      LAYER MET2 ;
        RECT 1.855 5.415 1.955 6 ;
      LAYER CUT12 ;
        RECT 1.855 5.765 1.955 5.865 ;
        RECT 1.855 5.545 1.955 5.645 ;
      LAYER CUT01 ;
        RECT 1.86 5.675 1.95 5.765 ;
        RECT 1.86 5.455 1.95 5.545 ;
    END
  END A
  PIN VDDSRC
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 3.79 3.79 5.23 11.57 ;
        RECT 3.79 3.79 11.57 5.23 ;
        RECT 2.2 2.2 3.64 11.57 ;
        RECT 2.2 2.2 11.57 3.64 ;
      LAYER CUT12 ;
        RECT 2.32 7.26 2.42 7.36 ;
        RECT 2.32 7.04 2.42 7.14 ;
        RECT 2.54 7.26 2.64 7.36 ;
        RECT 2.54 7.04 2.64 7.14 ;
        RECT 2.76 7.26 2.86 7.36 ;
        RECT 2.76 7.04 2.86 7.14 ;
        RECT 2.98 7.26 3.08 7.36 ;
        RECT 2.98 7.04 3.08 7.14 ;
        RECT 3.2 7.26 3.3 7.36 ;
        RECT 3.2 7.04 3.3 7.14 ;
        RECT 3.42 7.26 3.52 7.36 ;
        RECT 3.42 7.04 3.52 7.14 ;
        RECT 3.91 7.26 4.01 7.36 ;
        RECT 3.91 7.04 4.01 7.14 ;
        RECT 4.13 7.26 4.23 7.36 ;
        RECT 4.13 7.04 4.23 7.14 ;
        RECT 4.35 7.26 4.45 7.36 ;
        RECT 4.35 7.04 4.45 7.14 ;
        RECT 4.57 7.26 4.67 7.36 ;
        RECT 4.57 7.04 4.67 7.14 ;
        RECT 4.79 7.26 4.89 7.36 ;
        RECT 4.79 7.04 4.89 7.14 ;
        RECT 5.01 7.26 5.11 7.36 ;
        RECT 5.01 7.04 5.11 7.14 ;
        RECT 5.74 5.09 5.84 5.19 ;
        RECT 5.74 4.87 5.84 4.97 ;
        RECT 5.74 4.65 5.84 4.75 ;
        RECT 5.74 4.43 5.84 4.53 ;
    END
  END VDDSRC
  PIN Y
    DIRECTION OUTPUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNADIFFAREA 0.048 LAYER MET2 ;
    PORT
      LAYER MET1 ;
        RECT 5.47 5.43 5.57 10.89 ;
      LAYER MET2 ;
        RECT 5.38 5.38 6.48 11.57 ;
        RECT 5.38 5.38 11.57 6.48 ;
      LAYER CUT12 ;
        RECT 5.47 10.75 5.57 10.85 ;
        RECT 5.47 10.53 5.57 10.63 ;
        RECT 5.47 10.31 5.57 10.41 ;
        RECT 5.47 10.09 5.57 10.19 ;
        RECT 5.47 9.87 5.57 9.97 ;
        RECT 5.47 9.65 5.57 9.75 ;
        RECT 5.47 9.43 5.57 9.53 ;
        RECT 5.47 9.21 5.57 9.31 ;
        RECT 5.47 8.99 5.57 9.09 ;
        RECT 5.47 8.77 5.57 8.87 ;
        RECT 5.47 8.55 5.57 8.65 ;
        RECT 5.47 8.33 5.57 8.43 ;
        RECT 5.47 8.11 5.57 8.21 ;
        RECT 5.47 7.89 5.57 7.99 ;
        RECT 5.47 7.67 5.57 7.77 ;
        RECT 5.47 7.45 5.57 7.55 ;
        RECT 5.47 7.23 5.57 7.33 ;
        RECT 5.47 7.01 5.57 7.11 ;
        RECT 5.47 6.79 5.57 6.89 ;
        RECT 5.47 6.57 5.57 6.67 ;
        RECT 5.47 6.35 5.57 6.45 ;
        RECT 5.47 6.13 5.57 6.23 ;
        RECT 5.47 5.91 5.57 6.01 ;
        RECT 5.47 5.69 5.57 5.79 ;
        RECT 5.47 5.47 5.57 5.57 ;
      LAYER CUT01 ;
        RECT 5.475 6.375 5.565 6.465 ;
        RECT 5.475 5.605 5.565 5.695 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.28 0.37 2.38 5.71 ;
      RECT 1.855 5.415 1.955 6 ;
      RECT 1.855 5.9 2.44 6 ;
      RECT 2.34 5.865 2.44 6.035 ;
      RECT 2.28 6.41 2.38 7.36 ;
      RECT 2.28 7.04 5.15 7.36 ;
      RECT 2.55 5.9 5.37 6 ;
      RECT 5.27 5.865 5.37 6.035 ;
      RECT 2.55 5.59 2.65 6.42 ;
      RECT 5.47 5.43 5.57 10.89 ;
      RECT 5.74 5.88 6.46 5.98 ;
      RECT 5.74 4.39 5.84 6.505 ;
      RECT 6.54 0.37 6.64 5.71 ;
  END
END DSIPGX2LBFC1
MACRO DSIPGX2LBFF1
  CLASS RING ;
  ORIGIN 0 0 ;
  FOREIGN DSIPGX2LBFF1 0 0 ;
  SIZE 11.57 BY 11.57 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.23 0.23 0.37 11.57 ;
        RECT 0.23 0.23 11.57 0.37 ;
      LAYER CUT01 ;
        RECT 0.255 11.255 0.345 11.345 ;
        RECT 0.255 11.035 0.345 11.125 ;
        RECT 0.255 10.815 0.345 10.905 ;
        RECT 0.255 10.595 0.345 10.685 ;
        RECT 0.255 10.375 0.345 10.465 ;
        RECT 0.255 10.155 0.345 10.245 ;
        RECT 0.255 9.935 0.345 10.025 ;
        RECT 0.255 9.715 0.345 9.805 ;
        RECT 0.255 9.495 0.345 9.585 ;
        RECT 0.255 9.275 0.345 9.365 ;
        RECT 0.255 9.055 0.345 9.145 ;
        RECT 0.255 8.835 0.345 8.925 ;
        RECT 0.255 8.615 0.345 8.705 ;
        RECT 0.255 8.395 0.345 8.485 ;
        RECT 0.255 8.175 0.345 8.265 ;
        RECT 0.255 7.955 0.345 8.045 ;
        RECT 0.255 7.735 0.345 7.825 ;
        RECT 0.255 7.515 0.345 7.605 ;
        RECT 0.255 7.295 0.345 7.385 ;
        RECT 0.255 7.075 0.345 7.165 ;
        RECT 0.255 6.855 0.345 6.945 ;
        RECT 0.255 6.635 0.345 6.725 ;
        RECT 0.255 6.415 0.345 6.505 ;
        RECT 0.255 6.195 0.345 6.285 ;
        RECT 0.255 5.975 0.345 6.065 ;
        RECT 0.255 5.755 0.345 5.845 ;
        RECT 0.255 5.535 0.345 5.625 ;
        RECT 0.255 5.315 0.345 5.405 ;
        RECT 0.255 5.095 0.345 5.185 ;
        RECT 0.255 4.875 0.345 4.965 ;
        RECT 0.255 4.655 0.345 4.745 ;
        RECT 0.255 4.435 0.345 4.525 ;
        RECT 0.255 4.215 0.345 4.305 ;
        RECT 0.255 3.995 0.345 4.085 ;
        RECT 0.255 3.775 0.345 3.865 ;
        RECT 0.255 3.555 0.345 3.645 ;
        RECT 0.255 3.335 0.345 3.425 ;
        RECT 0.255 3.115 0.345 3.205 ;
        RECT 0.255 2.895 0.345 2.985 ;
        RECT 0.255 2.675 0.345 2.765 ;
        RECT 0.255 2.455 0.345 2.545 ;
        RECT 0.255 2.235 0.345 2.325 ;
        RECT 0.255 2.015 0.345 2.105 ;
        RECT 0.255 1.795 0.345 1.885 ;
        RECT 0.255 1.575 0.345 1.665 ;
        RECT 0.255 1.355 0.345 1.445 ;
        RECT 0.255 1.135 0.345 1.225 ;
        RECT 0.255 0.915 0.345 1.005 ;
        RECT 0.255 0.695 0.345 0.785 ;
        RECT 0.255 0.475 0.345 0.565 ;
        RECT 0.475 0.255 0.565 0.345 ;
        RECT 0.695 0.255 0.785 0.345 ;
        RECT 0.915 0.255 1.005 0.345 ;
        RECT 1.135 0.255 1.225 0.345 ;
        RECT 1.355 0.255 1.445 0.345 ;
        RECT 1.575 0.255 1.665 0.345 ;
        RECT 1.795 0.255 1.885 0.345 ;
        RECT 2.015 0.255 2.105 0.345 ;
        RECT 2.235 0.255 2.325 0.345 ;
        RECT 2.455 0.255 2.545 0.345 ;
        RECT 2.675 0.255 2.765 0.345 ;
        RECT 2.895 0.255 2.985 0.345 ;
        RECT 3.115 0.255 3.205 0.345 ;
        RECT 3.335 0.255 3.425 0.345 ;
        RECT 3.555 0.255 3.645 0.345 ;
        RECT 3.775 0.255 3.865 0.345 ;
        RECT 3.995 0.255 4.085 0.345 ;
        RECT 4.215 0.255 4.305 0.345 ;
        RECT 4.435 0.255 4.525 0.345 ;
        RECT 4.655 0.255 4.745 0.345 ;
        RECT 4.875 0.255 4.965 0.345 ;
        RECT 5.095 0.255 5.185 0.345 ;
        RECT 5.315 0.255 5.405 0.345 ;
        RECT 5.535 0.255 5.625 0.345 ;
        RECT 5.755 0.255 5.845 0.345 ;
        RECT 5.975 0.255 6.065 0.345 ;
        RECT 6.195 0.255 6.285 0.345 ;
        RECT 6.415 0.255 6.505 0.345 ;
        RECT 6.635 0.255 6.725 0.345 ;
        RECT 6.855 0.255 6.945 0.345 ;
        RECT 7.075 0.255 7.165 0.345 ;
        RECT 7.295 0.255 7.385 0.345 ;
        RECT 7.515 0.255 7.605 0.345 ;
        RECT 7.735 0.255 7.825 0.345 ;
        RECT 7.955 0.255 8.045 0.345 ;
        RECT 8.175 0.255 8.265 0.345 ;
        RECT 8.395 0.255 8.485 0.345 ;
        RECT 8.615 0.255 8.705 0.345 ;
        RECT 8.835 0.255 8.925 0.345 ;
        RECT 9.055 0.255 9.145 0.345 ;
        RECT 9.275 0.255 9.365 0.345 ;
        RECT 9.495 0.255 9.585 0.345 ;
        RECT 9.715 0.255 9.805 0.345 ;
        RECT 9.935 0.255 10.025 0.345 ;
        RECT 10.155 0.255 10.245 0.345 ;
        RECT 10.375 0.255 10.465 0.345 ;
        RECT 10.595 0.255 10.685 0.345 ;
        RECT 10.815 0.255 10.905 0.345 ;
        RECT 11.035 0.255 11.125 0.345 ;
        RECT 11.255 0.255 11.345 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 0.036 LAYER MET1 ;
      ANTENNAGATEAREA 0.036 LAYER MET2 ;
    ANTENNAMAXCUTCAR 416.666667 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDDSRC ;
    PORT
      LAYER MET1 ;
        RECT 1.855 5.415 1.955 6 ;
        RECT 1.855 5.9 2.44 6 ;
        RECT 2.34 5.865 2.44 6.035 ;
      LAYER MET2 ;
        RECT 1.855 5.415 1.955 6 ;
      LAYER CUT12 ;
        RECT 1.855 5.765 1.955 5.865 ;
        RECT 1.855 5.545 1.955 5.645 ;
      LAYER CUT01 ;
        RECT 1.86 5.675 1.95 5.765 ;
        RECT 1.86 5.455 1.95 5.545 ;
        RECT 2.345 5.905 2.435 5.995 ;
    END
  END A
  PIN VDDSRC
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 3.79 3.79 5.23 11.57 ;
        RECT 3.79 3.79 11.57 5.23 ;
        RECT 2.2 2.2 3.64 11.57 ;
        RECT 2.2 2.2 11.57 3.64 ;
      LAYER CUT12 ;
        RECT 2.32 7.26 2.42 7.36 ;
        RECT 2.32 7.04 2.42 7.14 ;
        RECT 2.54 7.26 2.64 7.36 ;
        RECT 2.54 7.04 2.64 7.14 ;
        RECT 2.76 7.26 2.86 7.36 ;
        RECT 2.76 7.04 2.86 7.14 ;
        RECT 2.98 7.26 3.08 7.36 ;
        RECT 2.98 7.04 3.08 7.14 ;
        RECT 3.2 7.26 3.3 7.36 ;
        RECT 3.2 7.04 3.3 7.14 ;
        RECT 3.42 7.26 3.52 7.36 ;
        RECT 3.42 7.04 3.52 7.14 ;
        RECT 3.91 7.26 4.01 7.36 ;
        RECT 3.91 7.04 4.01 7.14 ;
        RECT 4.13 7.26 4.23 7.36 ;
        RECT 4.13 7.04 4.23 7.14 ;
        RECT 4.35 7.26 4.45 7.36 ;
        RECT 4.35 7.04 4.45 7.14 ;
        RECT 4.57 7.26 4.67 7.36 ;
        RECT 4.57 7.04 4.67 7.14 ;
        RECT 4.79 7.26 4.89 7.36 ;
        RECT 4.79 7.04 4.89 7.14 ;
        RECT 5.01 7.26 5.11 7.36 ;
        RECT 5.01 7.04 5.11 7.14 ;
        RECT 5.74 5.09 5.84 5.19 ;
        RECT 5.74 4.87 5.84 4.97 ;
        RECT 5.74 4.65 5.84 4.75 ;
        RECT 5.74 4.43 5.84 4.53 ;
    END
  END VDDSRC
  PIN Y
    DIRECTION OUTPUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNADIFFAREA 0.048 LAYER MET2 ;
    PORT
      LAYER MET1 ;
        RECT 5.47 5.43 5.57 10.89 ;
      LAYER MET2 ;
        RECT 5.38 5.38 6.48 11.57 ;
        RECT 5.38 5.38 11.57 6.48 ;
      LAYER CUT12 ;
        RECT 5.47 10.75 5.57 10.85 ;
        RECT 5.47 10.53 5.57 10.63 ;
        RECT 5.47 10.31 5.57 10.41 ;
        RECT 5.47 10.09 5.57 10.19 ;
        RECT 5.47 9.87 5.57 9.97 ;
        RECT 5.47 9.65 5.57 9.75 ;
        RECT 5.47 9.43 5.57 9.53 ;
        RECT 5.47 9.21 5.57 9.31 ;
        RECT 5.47 8.99 5.57 9.09 ;
        RECT 5.47 8.77 5.57 8.87 ;
        RECT 5.47 8.55 5.57 8.65 ;
        RECT 5.47 8.33 5.57 8.43 ;
        RECT 5.47 8.11 5.57 8.21 ;
        RECT 5.47 7.89 5.57 7.99 ;
        RECT 5.47 7.67 5.57 7.77 ;
        RECT 5.47 7.45 5.57 7.55 ;
        RECT 5.47 7.23 5.57 7.33 ;
        RECT 5.47 7.01 5.57 7.11 ;
        RECT 5.47 6.79 5.57 6.89 ;
        RECT 5.47 6.57 5.57 6.67 ;
        RECT 5.47 6.35 5.57 6.45 ;
        RECT 5.47 6.13 5.57 6.23 ;
        RECT 5.47 5.91 5.57 6.01 ;
        RECT 5.47 5.69 5.57 5.79 ;
        RECT 5.47 5.47 5.57 5.57 ;
      LAYER CUT01 ;
        RECT 5.475 6.375 5.565 6.465 ;
        RECT 5.475 5.605 5.565 5.695 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.28 0.37 2.38 5.71 ;
      RECT 1.855 5.415 1.955 6 ;
      RECT 1.855 5.9 2.44 6 ;
      RECT 2.34 5.865 2.44 6.035 ;
      RECT 2.28 6.41 2.38 7.36 ;
      RECT 2.28 7.04 5.15 7.36 ;
      RECT 2.55 5.9 5.37 6 ;
      RECT 5.27 5.865 5.37 6.035 ;
      RECT 2.55 5.59 2.65 6.42 ;
      RECT 5.47 5.43 5.57 10.89 ;
      RECT 5.74 5.88 6.04 5.98 ;
      RECT 5.74 4.39 5.84 6.505 ;
      RECT 6.14 0.37 6.24 5.71 ;
  END
END DSIPGX2LBFF1
MACRO DSIPGX2LBFJ1
  CLASS RING ;
  ORIGIN 0 0 ;
  FOREIGN DSIPGX2LBFJ1 0 0 ;
  SIZE 11.57 BY 11.57 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.23 0.23 0.37 11.57 ;
        RECT 0.23 0.23 11.57 0.37 ;
      LAYER CUT01 ;
        RECT 0.255 11.255 0.345 11.345 ;
        RECT 0.255 11.035 0.345 11.125 ;
        RECT 0.255 10.815 0.345 10.905 ;
        RECT 0.255 10.595 0.345 10.685 ;
        RECT 0.255 10.375 0.345 10.465 ;
        RECT 0.255 10.155 0.345 10.245 ;
        RECT 0.255 9.935 0.345 10.025 ;
        RECT 0.255 9.715 0.345 9.805 ;
        RECT 0.255 9.495 0.345 9.585 ;
        RECT 0.255 9.275 0.345 9.365 ;
        RECT 0.255 9.055 0.345 9.145 ;
        RECT 0.255 8.835 0.345 8.925 ;
        RECT 0.255 8.615 0.345 8.705 ;
        RECT 0.255 8.395 0.345 8.485 ;
        RECT 0.255 8.175 0.345 8.265 ;
        RECT 0.255 7.955 0.345 8.045 ;
        RECT 0.255 7.735 0.345 7.825 ;
        RECT 0.255 7.515 0.345 7.605 ;
        RECT 0.255 7.295 0.345 7.385 ;
        RECT 0.255 7.075 0.345 7.165 ;
        RECT 0.255 6.855 0.345 6.945 ;
        RECT 0.255 6.635 0.345 6.725 ;
        RECT 0.255 6.415 0.345 6.505 ;
        RECT 0.255 6.195 0.345 6.285 ;
        RECT 0.255 5.975 0.345 6.065 ;
        RECT 0.255 5.755 0.345 5.845 ;
        RECT 0.255 5.535 0.345 5.625 ;
        RECT 0.255 5.315 0.345 5.405 ;
        RECT 0.255 5.095 0.345 5.185 ;
        RECT 0.255 4.875 0.345 4.965 ;
        RECT 0.255 4.655 0.345 4.745 ;
        RECT 0.255 4.435 0.345 4.525 ;
        RECT 0.255 4.215 0.345 4.305 ;
        RECT 0.255 3.995 0.345 4.085 ;
        RECT 0.255 3.775 0.345 3.865 ;
        RECT 0.255 3.555 0.345 3.645 ;
        RECT 0.255 3.335 0.345 3.425 ;
        RECT 0.255 3.115 0.345 3.205 ;
        RECT 0.255 2.895 0.345 2.985 ;
        RECT 0.255 2.675 0.345 2.765 ;
        RECT 0.255 2.455 0.345 2.545 ;
        RECT 0.255 2.235 0.345 2.325 ;
        RECT 0.255 2.015 0.345 2.105 ;
        RECT 0.255 1.795 0.345 1.885 ;
        RECT 0.255 1.575 0.345 1.665 ;
        RECT 0.255 1.355 0.345 1.445 ;
        RECT 0.255 1.135 0.345 1.225 ;
        RECT 0.255 0.915 0.345 1.005 ;
        RECT 0.255 0.695 0.345 0.785 ;
        RECT 0.255 0.475 0.345 0.565 ;
        RECT 0.475 0.255 0.565 0.345 ;
        RECT 0.695 0.255 0.785 0.345 ;
        RECT 0.915 0.255 1.005 0.345 ;
        RECT 1.135 0.255 1.225 0.345 ;
        RECT 1.355 0.255 1.445 0.345 ;
        RECT 1.575 0.255 1.665 0.345 ;
        RECT 1.795 0.255 1.885 0.345 ;
        RECT 2.015 0.255 2.105 0.345 ;
        RECT 2.235 0.255 2.325 0.345 ;
        RECT 2.455 0.255 2.545 0.345 ;
        RECT 2.675 0.255 2.765 0.345 ;
        RECT 2.895 0.255 2.985 0.345 ;
        RECT 3.115 0.255 3.205 0.345 ;
        RECT 3.335 0.255 3.425 0.345 ;
        RECT 3.555 0.255 3.645 0.345 ;
        RECT 3.775 0.255 3.865 0.345 ;
        RECT 3.995 0.255 4.085 0.345 ;
        RECT 4.215 0.255 4.305 0.345 ;
        RECT 4.435 0.255 4.525 0.345 ;
        RECT 4.655 0.255 4.745 0.345 ;
        RECT 4.875 0.255 4.965 0.345 ;
        RECT 5.095 0.255 5.185 0.345 ;
        RECT 5.315 0.255 5.405 0.345 ;
        RECT 5.535 0.255 5.625 0.345 ;
        RECT 5.755 0.255 5.845 0.345 ;
        RECT 5.975 0.255 6.065 0.345 ;
        RECT 6.195 0.255 6.285 0.345 ;
        RECT 6.415 0.255 6.505 0.345 ;
        RECT 6.635 0.255 6.725 0.345 ;
        RECT 6.855 0.255 6.945 0.345 ;
        RECT 7.075 0.255 7.165 0.345 ;
        RECT 7.295 0.255 7.385 0.345 ;
        RECT 7.515 0.255 7.605 0.345 ;
        RECT 7.735 0.255 7.825 0.345 ;
        RECT 7.955 0.255 8.045 0.345 ;
        RECT 8.175 0.255 8.265 0.345 ;
        RECT 8.395 0.255 8.485 0.345 ;
        RECT 8.615 0.255 8.705 0.345 ;
        RECT 8.835 0.255 8.925 0.345 ;
        RECT 9.055 0.255 9.145 0.345 ;
        RECT 9.275 0.255 9.365 0.345 ;
        RECT 9.495 0.255 9.585 0.345 ;
        RECT 9.715 0.255 9.805 0.345 ;
        RECT 9.935 0.255 10.025 0.345 ;
        RECT 10.155 0.255 10.245 0.345 ;
        RECT 10.375 0.255 10.465 0.345 ;
        RECT 10.595 0.255 10.685 0.345 ;
        RECT 10.815 0.255 10.905 0.345 ;
        RECT 11.035 0.255 11.125 0.345 ;
        RECT 11.255 0.255 11.345 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 0.036 LAYER MET1 ;
      ANTENNAGATEAREA 0.036 LAYER MET2 ;
    ANTENNAMAXCUTCAR 416.666667 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDDSRC ;
    PORT
      LAYER MET1 ;
        RECT 1.855 5.415 1.955 6 ;
        RECT 1.855 5.9 2.44 6 ;
        RECT 2.34 5.865 2.44 6.035 ;
      LAYER MET2 ;
        RECT 1.855 5.415 1.955 6 ;
      LAYER CUT12 ;
        RECT 1.855 5.765 1.955 5.865 ;
        RECT 1.855 5.545 1.955 5.645 ;
      LAYER CUT01 ;
        RECT 1.86 5.675 1.95 5.765 ;
        RECT 1.86 5.455 1.95 5.545 ;
        RECT 2.345 5.905 2.435 5.995 ;
    END
  END A
  PIN VDDSRC
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 3.79 3.79 5.23 11.57 ;
        RECT 3.79 3.79 11.57 5.23 ;
        RECT 2.2 2.2 3.64 11.57 ;
        RECT 2.2 2.2 11.57 3.64 ;
      LAYER CUT12 ;
        RECT 2.32 7.26 2.42 7.36 ;
        RECT 2.32 7.04 2.42 7.14 ;
        RECT 2.54 7.26 2.64 7.36 ;
        RECT 2.54 7.04 2.64 7.14 ;
        RECT 2.76 7.26 2.86 7.36 ;
        RECT 2.76 7.04 2.86 7.14 ;
        RECT 2.98 7.26 3.08 7.36 ;
        RECT 2.98 7.04 3.08 7.14 ;
        RECT 3.2 7.26 3.3 7.36 ;
        RECT 3.2 7.04 3.3 7.14 ;
        RECT 3.42 7.26 3.52 7.36 ;
        RECT 3.42 7.04 3.52 7.14 ;
        RECT 3.91 7.26 4.01 7.36 ;
        RECT 3.91 7.04 4.01 7.14 ;
        RECT 4.13 7.26 4.23 7.36 ;
        RECT 4.13 7.04 4.23 7.14 ;
        RECT 4.35 7.26 4.45 7.36 ;
        RECT 4.35 7.04 4.45 7.14 ;
        RECT 4.57 7.26 4.67 7.36 ;
        RECT 4.57 7.04 4.67 7.14 ;
        RECT 4.79 7.26 4.89 7.36 ;
        RECT 4.79 7.04 4.89 7.14 ;
        RECT 5.01 7.26 5.11 7.36 ;
        RECT 5.01 7.04 5.11 7.14 ;
        RECT 6.04 5.09 6.14 5.19 ;
        RECT 6.04 4.87 6.14 4.97 ;
        RECT 6.04 4.65 6.14 4.75 ;
        RECT 6.04 4.43 6.14 4.53 ;
    END
  END VDDSRC
  PIN Y
    DIRECTION OUTPUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 0.048 LAYER MET1 ;
    ANTENNADIFFAREA 0.048 LAYER MET2 ;
    PORT
      LAYER MET1 ;
        RECT 5.47 5.43 5.57 10.89 ;
      LAYER MET2 ;
        RECT 5.38 5.38 6.48 11.57 ;
        RECT 5.38 5.38 11.57 6.48 ;
      LAYER CUT12 ;
        RECT 5.47 10.75 5.57 10.85 ;
        RECT 5.47 10.53 5.57 10.63 ;
        RECT 5.47 10.31 5.57 10.41 ;
        RECT 5.47 10.09 5.57 10.19 ;
        RECT 5.47 9.87 5.57 9.97 ;
        RECT 5.47 9.65 5.57 9.75 ;
        RECT 5.47 9.43 5.57 9.53 ;
        RECT 5.47 9.21 5.57 9.31 ;
        RECT 5.47 8.99 5.57 9.09 ;
        RECT 5.47 8.77 5.57 8.87 ;
        RECT 5.47 8.55 5.57 8.65 ;
        RECT 5.47 8.33 5.57 8.43 ;
        RECT 5.47 8.11 5.57 8.21 ;
        RECT 5.47 7.89 5.57 7.99 ;
        RECT 5.47 7.67 5.57 7.77 ;
        RECT 5.47 7.45 5.57 7.55 ;
        RECT 5.47 7.23 5.57 7.33 ;
        RECT 5.47 7.01 5.57 7.11 ;
        RECT 5.47 6.79 5.57 6.89 ;
        RECT 5.47 6.57 5.57 6.67 ;
        RECT 5.47 6.35 5.57 6.45 ;
        RECT 5.47 6.13 5.57 6.23 ;
        RECT 5.47 5.91 5.57 6.01 ;
        RECT 5.47 5.69 5.57 5.79 ;
        RECT 5.47 5.47 5.57 5.57 ;
      LAYER CUT01 ;
        RECT 5.475 6.375 5.565 6.465 ;
        RECT 5.475 5.605 5.565 5.695 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.28 0.37 2.38 5.71 ;
      RECT 1.855 5.415 1.955 6 ;
      RECT 1.855 5.9 2.44 6 ;
      RECT 2.34 5.865 2.44 6.035 ;
      RECT 2.28 6.41 2.38 7.36 ;
      RECT 2.28 7.04 5.15 7.36 ;
      RECT 2.55 5.9 5.37 6 ;
      RECT 5.27 5.865 5.37 6.035 ;
      RECT 2.55 5.59 2.65 6.42 ;
      RECT 5.47 5.43 5.57 10.89 ;
      RECT 5.74 0.37 5.84 5.71 ;
      RECT 6.04 4.39 6.14 6 ;
      RECT 5.74 5.9 6.14 6 ;
      RECT 5.74 5.9 5.84 6.505 ;
  END
END DSIPGX2LBFJ1
MACRO DSIPGX2LBFL1
  CLASS RING ;
  ORIGIN 0 0 ;
  FOREIGN DSIPGX2LBFL1 0 0 ;
  SIZE 11.57 BY 11.57 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.23 0.23 0.37 11.57 ;
        RECT 0.23 0.23 11.57 0.37 ;
      LAYER CUT01 ;
        RECT 0.255 11.255 0.345 11.345 ;
        RECT 0.255 11.035 0.345 11.125 ;
        RECT 0.255 10.815 0.345 10.905 ;
        RECT 0.255 10.595 0.345 10.685 ;
        RECT 0.255 10.375 0.345 10.465 ;
        RECT 0.255 10.155 0.345 10.245 ;
        RECT 0.255 9.935 0.345 10.025 ;
        RECT 0.255 9.715 0.345 9.805 ;
        RECT 0.255 9.495 0.345 9.585 ;
        RECT 0.255 9.275 0.345 9.365 ;
        RECT 0.255 9.055 0.345 9.145 ;
        RECT 0.255 8.835 0.345 8.925 ;
        RECT 0.255 8.615 0.345 8.705 ;
        RECT 0.255 8.395 0.345 8.485 ;
        RECT 0.255 8.175 0.345 8.265 ;
        RECT 0.255 7.955 0.345 8.045 ;
        RECT 0.255 7.735 0.345 7.825 ;
        RECT 0.255 7.515 0.345 7.605 ;
        RECT 0.255 7.295 0.345 7.385 ;
        RECT 0.255 7.075 0.345 7.165 ;
        RECT 0.255 6.855 0.345 6.945 ;
        RECT 0.255 6.635 0.345 6.725 ;
        RECT 0.255 6.415 0.345 6.505 ;
        RECT 0.255 6.195 0.345 6.285 ;
        RECT 0.255 5.975 0.345 6.065 ;
        RECT 0.255 5.755 0.345 5.845 ;
        RECT 0.255 5.535 0.345 5.625 ;
        RECT 0.255 5.315 0.345 5.405 ;
        RECT 0.255 5.095 0.345 5.185 ;
        RECT 0.255 4.875 0.345 4.965 ;
        RECT 0.255 4.655 0.345 4.745 ;
        RECT 0.255 4.435 0.345 4.525 ;
        RECT 0.255 4.215 0.345 4.305 ;
        RECT 0.255 3.995 0.345 4.085 ;
        RECT 0.255 3.775 0.345 3.865 ;
        RECT 0.255 3.555 0.345 3.645 ;
        RECT 0.255 3.335 0.345 3.425 ;
        RECT 0.255 3.115 0.345 3.205 ;
        RECT 0.255 2.895 0.345 2.985 ;
        RECT 0.255 2.675 0.345 2.765 ;
        RECT 0.255 2.455 0.345 2.545 ;
        RECT 0.255 2.235 0.345 2.325 ;
        RECT 0.255 2.015 0.345 2.105 ;
        RECT 0.255 1.795 0.345 1.885 ;
        RECT 0.255 1.575 0.345 1.665 ;
        RECT 0.255 1.355 0.345 1.445 ;
        RECT 0.255 1.135 0.345 1.225 ;
        RECT 0.255 0.915 0.345 1.005 ;
        RECT 0.255 0.695 0.345 0.785 ;
        RECT 0.255 0.475 0.345 0.565 ;
        RECT 0.475 0.255 0.565 0.345 ;
        RECT 0.695 0.255 0.785 0.345 ;
        RECT 0.915 0.255 1.005 0.345 ;
        RECT 1.135 0.255 1.225 0.345 ;
        RECT 1.355 0.255 1.445 0.345 ;
        RECT 1.575 0.255 1.665 0.345 ;
        RECT 1.795 0.255 1.885 0.345 ;
        RECT 2.015 0.255 2.105 0.345 ;
        RECT 2.235 0.255 2.325 0.345 ;
        RECT 2.455 0.255 2.545 0.345 ;
        RECT 2.675 0.255 2.765 0.345 ;
        RECT 2.895 0.255 2.985 0.345 ;
        RECT 3.115 0.255 3.205 0.345 ;
        RECT 3.335 0.255 3.425 0.345 ;
        RECT 3.555 0.255 3.645 0.345 ;
        RECT 3.775 0.255 3.865 0.345 ;
        RECT 3.995 0.255 4.085 0.345 ;
        RECT 4.215 0.255 4.305 0.345 ;
        RECT 4.435 0.255 4.525 0.345 ;
        RECT 4.655 0.255 4.745 0.345 ;
        RECT 4.875 0.255 4.965 0.345 ;
        RECT 5.095 0.255 5.185 0.345 ;
        RECT 5.315 0.255 5.405 0.345 ;
        RECT 5.535 0.255 5.625 0.345 ;
        RECT 5.755 0.255 5.845 0.345 ;
        RECT 5.975 0.255 6.065 0.345 ;
        RECT 6.195 0.255 6.285 0.345 ;
        RECT 6.415 0.255 6.505 0.345 ;
        RECT 6.635 0.255 6.725 0.345 ;
        RECT 6.855 0.255 6.945 0.345 ;
        RECT 7.075 0.255 7.165 0.345 ;
        RECT 7.295 0.255 7.385 0.345 ;
        RECT 7.515 0.255 7.605 0.345 ;
        RECT 7.735 0.255 7.825 0.345 ;
        RECT 7.955 0.255 8.045 0.345 ;
        RECT 8.175 0.255 8.265 0.345 ;
        RECT 8.395 0.255 8.485 0.345 ;
        RECT 8.615 0.255 8.705 0.345 ;
        RECT 8.835 0.255 8.925 0.345 ;
        RECT 9.055 0.255 9.145 0.345 ;
        RECT 9.275 0.255 9.365 0.345 ;
        RECT 9.495 0.255 9.585 0.345 ;
        RECT 9.715 0.255 9.805 0.345 ;
        RECT 9.935 0.255 10.025 0.345 ;
        RECT 10.155 0.255 10.245 0.345 ;
        RECT 10.375 0.255 10.465 0.345 ;
        RECT 10.595 0.255 10.685 0.345 ;
        RECT 10.815 0.255 10.905 0.345 ;
        RECT 11.035 0.255 11.125 0.345 ;
        RECT 11.255 0.255 11.345 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 0.036 LAYER MET1 ;
      ANTENNAGATEAREA 0.036 LAYER MET2 ;
    ANTENNAMAXCUTCAR 416.666667 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDDSRC ;
    PORT
      LAYER MET1 ;
        RECT 1.855 5.415 1.955 6 ;
        RECT 1.855 5.9 2.44 6 ;
        RECT 2.34 5.865 2.44 6.035 ;
      LAYER MET2 ;
        RECT 1.855 5.415 1.955 6 ;
      LAYER CUT12 ;
        RECT 1.855 5.765 1.955 5.865 ;
        RECT 1.855 5.545 1.955 5.645 ;
      LAYER CUT01 ;
        RECT 1.86 5.675 1.95 5.765 ;
        RECT 1.86 5.455 1.95 5.545 ;
        RECT 2.345 5.905 2.435 5.995 ;
    END
  END A
  PIN VDDSRC
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 3.79 3.79 5.23 11.57 ;
        RECT 3.79 3.79 11.57 5.23 ;
        RECT 2.2 2.2 3.64 11.57 ;
        RECT 2.2 2.2 11.57 3.64 ;
      LAYER CUT12 ;
        RECT 2.32 7.26 2.42 7.36 ;
        RECT 2.32 7.04 2.42 7.14 ;
        RECT 2.54 7.26 2.64 7.36 ;
        RECT 2.54 7.04 2.64 7.14 ;
        RECT 2.76 7.26 2.86 7.36 ;
        RECT 2.76 7.04 2.86 7.14 ;
        RECT 2.98 7.26 3.08 7.36 ;
        RECT 2.98 7.04 3.08 7.14 ;
        RECT 3.2 7.26 3.3 7.36 ;
        RECT 3.2 7.04 3.3 7.14 ;
        RECT 3.42 7.26 3.52 7.36 ;
        RECT 3.42 7.04 3.52 7.14 ;
        RECT 3.91 7.26 4.01 7.36 ;
        RECT 3.91 7.04 4.01 7.14 ;
        RECT 4.13 7.26 4.23 7.36 ;
        RECT 4.13 7.04 4.23 7.14 ;
        RECT 4.35 7.26 4.45 7.36 ;
        RECT 4.35 7.04 4.45 7.14 ;
        RECT 4.57 7.26 4.67 7.36 ;
        RECT 4.57 7.04 4.67 7.14 ;
        RECT 4.79 7.26 4.89 7.36 ;
        RECT 4.79 7.04 4.89 7.14 ;
        RECT 5.01 7.26 5.11 7.36 ;
        RECT 5.01 7.04 5.11 7.14 ;
        RECT 6.04 5.09 6.14 5.19 ;
        RECT 6.04 4.87 6.14 4.97 ;
        RECT 6.04 4.65 6.14 4.75 ;
        RECT 6.04 4.43 6.14 4.53 ;
    END
  END VDDSRC
  PIN Y
    DIRECTION OUTPUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 0.0744 LAYER MET1 ;
    ANTENNADIFFAREA 0.0744 LAYER MET2 ;
    PORT
      LAYER MET1 ;
        RECT 5.47 5.37 5.57 10.89 ;
      LAYER MET2 ;
        RECT 5.38 5.38 6.48 11.57 ;
        RECT 5.38 5.38 11.57 6.48 ;
      LAYER CUT12 ;
        RECT 5.47 10.75 5.57 10.85 ;
        RECT 5.47 10.53 5.57 10.63 ;
        RECT 5.47 10.31 5.57 10.41 ;
        RECT 5.47 10.09 5.57 10.19 ;
        RECT 5.47 9.87 5.57 9.97 ;
        RECT 5.47 9.65 5.57 9.75 ;
        RECT 5.47 9.43 5.57 9.53 ;
        RECT 5.47 9.21 5.57 9.31 ;
        RECT 5.47 8.99 5.57 9.09 ;
        RECT 5.47 8.77 5.57 8.87 ;
        RECT 5.47 8.55 5.57 8.65 ;
        RECT 5.47 8.33 5.57 8.43 ;
        RECT 5.47 8.11 5.57 8.21 ;
        RECT 5.47 7.89 5.57 7.99 ;
        RECT 5.47 7.67 5.57 7.77 ;
        RECT 5.47 7.45 5.57 7.55 ;
        RECT 5.47 7.23 5.57 7.33 ;
        RECT 5.47 7.01 5.57 7.11 ;
        RECT 5.47 6.79 5.57 6.89 ;
        RECT 5.47 6.57 5.57 6.67 ;
        RECT 5.47 6.35 5.57 6.45 ;
        RECT 5.47 6.13 5.57 6.23 ;
        RECT 5.47 5.91 5.57 6.01 ;
        RECT 5.47 5.69 5.57 5.79 ;
        RECT 5.47 5.47 5.57 5.57 ;
      LAYER CUT01 ;
        RECT 5.475 6.625 5.565 6.715 ;
        RECT 5.475 6.405 5.565 6.495 ;
        RECT 5.475 6.185 5.565 6.275 ;
        RECT 5.475 5.63 5.565 5.72 ;
        RECT 5.475 5.41 5.565 5.5 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.28 0.37 2.38 5.71 ;
      RECT 1.855 5.415 1.955 6 ;
      RECT 1.855 5.9 2.44 6 ;
      RECT 2.34 5.865 2.44 6.035 ;
      RECT 2.28 6.41 2.38 7.36 ;
      RECT 2.28 7.04 5.15 7.36 ;
      RECT 2.55 5.9 5.37 6 ;
      RECT 5.27 5.865 5.37 6.035 ;
      RECT 2.55 5.59 2.65 6.42 ;
      RECT 5.47 5.37 5.57 10.89 ;
      RECT 5.74 0.37 5.84 5.76 ;
      RECT 6.04 4.39 6.14 6 ;
      RECT 5.74 5.9 6.14 6 ;
      RECT 5.74 5.9 5.84 6.755 ;
  END
END DSIPGX2LBFL1
MACRO DSIPGX2LBFN1
  CLASS RING ;
  ORIGIN 0 0 ;
  FOREIGN DSIPGX2LBFN1 0 0 ;
  SIZE 11.57 BY 11.57 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.23 0.23 0.37 11.57 ;
        RECT 0.23 0.23 11.57 0.37 ;
      LAYER CUT01 ;
        RECT 0.255 11.255 0.345 11.345 ;
        RECT 0.255 11.035 0.345 11.125 ;
        RECT 0.255 10.815 0.345 10.905 ;
        RECT 0.255 10.595 0.345 10.685 ;
        RECT 0.255 10.375 0.345 10.465 ;
        RECT 0.255 10.155 0.345 10.245 ;
        RECT 0.255 9.935 0.345 10.025 ;
        RECT 0.255 9.715 0.345 9.805 ;
        RECT 0.255 9.495 0.345 9.585 ;
        RECT 0.255 9.275 0.345 9.365 ;
        RECT 0.255 9.055 0.345 9.145 ;
        RECT 0.255 8.835 0.345 8.925 ;
        RECT 0.255 8.615 0.345 8.705 ;
        RECT 0.255 8.395 0.345 8.485 ;
        RECT 0.255 8.175 0.345 8.265 ;
        RECT 0.255 7.955 0.345 8.045 ;
        RECT 0.255 7.735 0.345 7.825 ;
        RECT 0.255 7.515 0.345 7.605 ;
        RECT 0.255 7.295 0.345 7.385 ;
        RECT 0.255 7.075 0.345 7.165 ;
        RECT 0.255 6.855 0.345 6.945 ;
        RECT 0.255 6.635 0.345 6.725 ;
        RECT 0.255 6.415 0.345 6.505 ;
        RECT 0.255 6.195 0.345 6.285 ;
        RECT 0.255 5.975 0.345 6.065 ;
        RECT 0.255 5.755 0.345 5.845 ;
        RECT 0.255 5.535 0.345 5.625 ;
        RECT 0.255 5.315 0.345 5.405 ;
        RECT 0.255 5.095 0.345 5.185 ;
        RECT 0.255 4.875 0.345 4.965 ;
        RECT 0.255 4.655 0.345 4.745 ;
        RECT 0.255 4.435 0.345 4.525 ;
        RECT 0.255 4.215 0.345 4.305 ;
        RECT 0.255 3.995 0.345 4.085 ;
        RECT 0.255 3.775 0.345 3.865 ;
        RECT 0.255 3.555 0.345 3.645 ;
        RECT 0.255 3.335 0.345 3.425 ;
        RECT 0.255 3.115 0.345 3.205 ;
        RECT 0.255 2.895 0.345 2.985 ;
        RECT 0.255 2.675 0.345 2.765 ;
        RECT 0.255 2.455 0.345 2.545 ;
        RECT 0.255 2.235 0.345 2.325 ;
        RECT 0.255 2.015 0.345 2.105 ;
        RECT 0.255 1.795 0.345 1.885 ;
        RECT 0.255 1.575 0.345 1.665 ;
        RECT 0.255 1.355 0.345 1.445 ;
        RECT 0.255 1.135 0.345 1.225 ;
        RECT 0.255 0.915 0.345 1.005 ;
        RECT 0.255 0.695 0.345 0.785 ;
        RECT 0.255 0.475 0.345 0.565 ;
        RECT 0.475 0.255 0.565 0.345 ;
        RECT 0.695 0.255 0.785 0.345 ;
        RECT 0.915 0.255 1.005 0.345 ;
        RECT 1.135 0.255 1.225 0.345 ;
        RECT 1.355 0.255 1.445 0.345 ;
        RECT 1.575 0.255 1.665 0.345 ;
        RECT 1.795 0.255 1.885 0.345 ;
        RECT 2.015 0.255 2.105 0.345 ;
        RECT 2.235 0.255 2.325 0.345 ;
        RECT 2.455 0.255 2.545 0.345 ;
        RECT 2.675 0.255 2.765 0.345 ;
        RECT 2.895 0.255 2.985 0.345 ;
        RECT 3.115 0.255 3.205 0.345 ;
        RECT 3.335 0.255 3.425 0.345 ;
        RECT 3.555 0.255 3.645 0.345 ;
        RECT 3.775 0.255 3.865 0.345 ;
        RECT 3.995 0.255 4.085 0.345 ;
        RECT 4.215 0.255 4.305 0.345 ;
        RECT 4.435 0.255 4.525 0.345 ;
        RECT 4.655 0.255 4.745 0.345 ;
        RECT 4.875 0.255 4.965 0.345 ;
        RECT 5.095 0.255 5.185 0.345 ;
        RECT 5.315 0.255 5.405 0.345 ;
        RECT 5.535 0.255 5.625 0.345 ;
        RECT 5.755 0.255 5.845 0.345 ;
        RECT 5.975 0.255 6.065 0.345 ;
        RECT 6.195 0.255 6.285 0.345 ;
        RECT 6.415 0.255 6.505 0.345 ;
        RECT 6.635 0.255 6.725 0.345 ;
        RECT 6.855 0.255 6.945 0.345 ;
        RECT 7.075 0.255 7.165 0.345 ;
        RECT 7.295 0.255 7.385 0.345 ;
        RECT 7.515 0.255 7.605 0.345 ;
        RECT 7.735 0.255 7.825 0.345 ;
        RECT 7.955 0.255 8.045 0.345 ;
        RECT 8.175 0.255 8.265 0.345 ;
        RECT 8.395 0.255 8.485 0.345 ;
        RECT 8.615 0.255 8.705 0.345 ;
        RECT 8.835 0.255 8.925 0.345 ;
        RECT 9.055 0.255 9.145 0.345 ;
        RECT 9.275 0.255 9.365 0.345 ;
        RECT 9.495 0.255 9.585 0.345 ;
        RECT 9.715 0.255 9.805 0.345 ;
        RECT 9.935 0.255 10.025 0.345 ;
        RECT 10.155 0.255 10.245 0.345 ;
        RECT 10.375 0.255 10.465 0.345 ;
        RECT 10.595 0.255 10.685 0.345 ;
        RECT 10.815 0.255 10.905 0.345 ;
        RECT 11.035 0.255 11.125 0.345 ;
        RECT 11.255 0.255 11.345 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
      ANTENNAGATEAREA 0.0507 LAYER MET1 ;
      ANTENNAGATEAREA 0.0507 LAYER MET2 ;
    ANTENNAMAXCUTCAR 295.857988 LAYER CUT01 ;
    GROUNDSENSITIVITY VSS ;
    SUPPLYSENSITIVITY VDDSRC ;
    PORT
      LAYER CUT01 ;
        RECT 2.345 5.905 2.435 5.995 ;
      LAYER MET1 ;
        RECT 1.855 5.415 1.955 6 ;
        RECT 1.855 5.9 2.44 6 ;
        RECT 2.34 5.865 2.44 6.035 ;
      LAYER MET2 ;
        RECT 1.855 5.415 1.955 6 ;
      LAYER CUT12 ;
        RECT 1.855 5.765 1.955 5.865 ;
        RECT 1.855 5.545 1.955 5.645 ;
      LAYER CUT01 ;
        RECT 1.86 5.675 1.95 5.765 ;
        RECT 1.86 5.455 1.95 5.545 ;
    END
  END A
  PIN VDDSRC
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 3.79 3.79 5.23 11.57 ;
        RECT 3.79 3.79 11.57 5.23 ;
        RECT 2.2 2.2 3.64 11.57 ;
        RECT 2.2 2.2 11.57 3.64 ;
      LAYER CUT12 ;
        RECT 2.32 7.26 2.42 7.36 ;
        RECT 2.32 7.04 2.42 7.14 ;
        RECT 2.54 7.26 2.64 7.36 ;
        RECT 2.54 7.04 2.64 7.14 ;
        RECT 2.76 7.26 2.86 7.36 ;
        RECT 2.76 7.04 2.86 7.14 ;
        RECT 2.98 7.26 3.08 7.36 ;
        RECT 2.98 7.04 3.08 7.14 ;
        RECT 3.2 7.26 3.3 7.36 ;
        RECT 3.2 7.04 3.3 7.14 ;
        RECT 3.42 7.26 3.52 7.36 ;
        RECT 3.42 7.04 3.52 7.14 ;
        RECT 3.91 7.26 4.01 7.36 ;
        RECT 3.91 7.04 4.01 7.14 ;
        RECT 4.13 7.26 4.23 7.36 ;
        RECT 4.13 7.04 4.23 7.14 ;
        RECT 4.35 7.26 4.45 7.36 ;
        RECT 4.35 7.04 4.45 7.14 ;
        RECT 4.57 7.26 4.67 7.36 ;
        RECT 4.57 7.04 4.67 7.14 ;
        RECT 4.79 7.26 4.89 7.36 ;
        RECT 4.79 7.04 4.89 7.14 ;
        RECT 5.01 7.26 5.11 7.36 ;
        RECT 5.01 7.04 5.11 7.14 ;
        RECT 6.04 5.09 6.14 5.19 ;
        RECT 6.04 4.87 6.14 4.97 ;
        RECT 6.04 4.65 6.14 4.75 ;
        RECT 6.04 4.43 6.14 4.53 ;
    END
  END VDDSRC
  PIN Y
    DIRECTION OUTPUT ;
    USE ANALOG ;
    ANTENNADIFFAREA 0.093 LAYER MET1 ;
    ANTENNADIFFAREA 0.093 LAYER MET2 ;
    PORT
      LAYER MET1 ;
        RECT 5.47 5.37 5.57 10.89 ;
      LAYER MET2 ;
        RECT 5.38 5.38 6.48 11.57 ;
        RECT 5.38 5.38 11.57 6.48 ;
      LAYER CUT12 ;
        RECT 5.47 10.75 5.57 10.85 ;
        RECT 5.47 10.53 5.57 10.63 ;
        RECT 5.47 10.31 5.57 10.41 ;
        RECT 5.47 10.09 5.57 10.19 ;
        RECT 5.47 9.87 5.57 9.97 ;
        RECT 5.47 9.65 5.57 9.75 ;
        RECT 5.47 9.43 5.57 9.53 ;
        RECT 5.47 9.21 5.57 9.31 ;
        RECT 5.47 8.99 5.57 9.09 ;
        RECT 5.47 8.77 5.57 8.87 ;
        RECT 5.47 8.55 5.57 8.65 ;
        RECT 5.47 8.33 5.57 8.43 ;
        RECT 5.47 8.11 5.57 8.21 ;
        RECT 5.47 7.89 5.57 7.99 ;
        RECT 5.47 7.67 5.57 7.77 ;
        RECT 5.47 7.45 5.57 7.55 ;
        RECT 5.47 7.23 5.57 7.33 ;
        RECT 5.47 7.01 5.57 7.11 ;
        RECT 5.47 6.79 5.57 6.89 ;
        RECT 5.47 6.57 5.57 6.67 ;
        RECT 5.47 6.35 5.57 6.45 ;
        RECT 5.47 6.13 5.57 6.23 ;
        RECT 5.47 5.91 5.57 6.01 ;
        RECT 5.47 5.69 5.57 5.79 ;
        RECT 5.47 5.47 5.57 5.57 ;
      LAYER CUT01 ;
        RECT 5.475 6.625 5.565 6.715 ;
        RECT 5.475 6.405 5.565 6.495 ;
        RECT 5.475 6.185 5.565 6.275 ;
        RECT 5.475 5.63 5.565 5.72 ;
        RECT 5.475 5.41 5.565 5.5 ;
    END
  END Y
  OBS
    LAYER MET1 ;
      RECT 2.28 0.37 2.38 5.685 ;
      RECT 1.855 5.415 1.955 6 ;
      RECT 1.855 5.9 2.44 6 ;
      RECT 2.34 5.865 2.44 6.035 ;
      RECT 2.28 6.3 2.38 7.36 ;
      RECT 5.2 6.145 5.3 7.36 ;
      RECT 2.28 7.04 5.3 7.36 ;
      RECT 2.55 5.9 5.37 6 ;
      RECT 5.27 5.865 5.37 6.035 ;
      RECT 2.55 5.515 2.65 6.69 ;
      RECT 5.47 5.37 5.57 10.89 ;
      RECT 5.2 4.905 5.84 5.005 ;
      RECT 5.2 4.905 5.3 5.76 ;
      RECT 5.74 0.37 5.84 5.76 ;
      RECT 6.04 4.39 6.14 6 ;
      RECT 5.74 5.9 6.14 6 ;
      RECT 5.74 5.9 5.84 6.755 ;
  END
END DSIPGX2LBFN1

MACRO DSIPGX2LPSCCS1
  CLASS CORE ;
  ORIGIN 0 0 ;
  FOREIGN DSIPGX2LPSCCS1 0 0 ;
  SIZE 9.8 BY 3.6 ;
  SYMMETRY X Y ;
  SITE WCORE3600 ;
  PIN A
    DIRECTION INPUT ;
    USE ANALOG ;
      ANTENNAGATEAREA 7.424 LAYER MET1 ;
    ANTENNAMAXCUTCAR 10.102371 LAYER CUT01 ;
    SUPPLYSENSITIVITY VDDSRC ;
    GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 0.08 3.19 9.72 3.29 ;
      LAYER CUT01 ;
        RECT 2.075 3.195 2.165 3.285 ;
        RECT 2.295 3.195 2.385 3.285 ;
        RECT 2.515 3.195 2.605 3.285 ;
        RECT 2.735 3.195 2.825 3.285 ;
        RECT 2.955 3.195 3.045 3.285 ;
        RECT 3.175 3.195 3.265 3.285 ;
        RECT 3.395 3.195 3.485 3.285 ;
        RECT 3.615 3.195 3.705 3.285 ;
        RECT 3.835 3.195 3.925 3.285 ;
        RECT 4.055 3.195 4.145 3.285 ;
        RECT 4.275 3.195 4.365 3.285 ;
        RECT 4.495 3.195 4.585 3.285 ;
        RECT 4.715 3.195 4.805 3.285 ;
        RECT 4.935 3.195 5.025 3.285 ;
        RECT 5.155 3.195 5.245 3.285 ;
        RECT 5.375 3.195 5.465 3.285 ;
        RECT 5.595 3.195 5.685 3.285 ;
        RECT 5.815 3.195 5.905 3.285 ;
        RECT 6.035 3.195 6.125 3.285 ;
        RECT 6.255 3.195 6.345 3.285 ;
        RECT 6.475 3.195 6.565 3.285 ;
        RECT 6.695 3.195 6.785 3.285 ;
        RECT 6.915 3.195 7.005 3.285 ;
        RECT 7.135 3.195 7.225 3.285 ;
        RECT 7.355 3.195 7.445 3.285 ;
    END
  END A
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 3.44 9.8 3.76 ;
        RECT 0 -0.16 9.8 0.16 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER CUT12 ;
        RECT 7.3 1.075 7.4 1.175 ;
        RECT 7.49 1.845 7.59 1.945 ;
        RECT 7.71 1.845 7.81 1.945 ;
        RECT 7.93 1.845 8.03 1.945 ;
        RECT 8.15 1.845 8.25 1.945 ;
        RECT 8.37 1.845 8.47 1.945 ;
        RECT 8.59 1.845 8.69 1.945 ;
        RECT 8.81 1.845 8.91 1.945 ;
        RECT 9.03 1.845 9.13 1.945 ;
        RECT 9.25 1.845 9.35 1.945 ;
        RECT 9.47 1.845 9.57 1.945 ;
      LAYER MET2 ;
        RECT 0.08 1.06 9.72 2.26 ;
      LAYER MET1 ;
        RECT 0 1.64 9.8 1.96 ;
      LAYER CUT01 ;
        RECT 2.125 1.905 2.215 1.995 ;
        RECT 2.125 1.685 2.215 1.775 ;
        RECT 2.865 1.905 2.955 1.995 ;
        RECT 2.865 1.685 2.955 1.775 ;
        RECT 3.605 1.905 3.695 1.995 ;
        RECT 3.605 1.685 3.695 1.775 ;
        RECT 4.345 1.905 4.435 1.995 ;
        RECT 4.345 1.685 4.435 1.775 ;
        RECT 5.085 1.905 5.175 1.995 ;
        RECT 5.085 1.685 5.175 1.775 ;
        RECT 5.825 1.905 5.915 1.995 ;
        RECT 5.825 1.685 5.915 1.775 ;
        RECT 6.565 1.905 6.655 1.995 ;
        RECT 6.565 1.685 6.655 1.775 ;
        RECT 7.305 1.905 7.395 1.995 ;
        RECT 7.305 1.685 7.395 1.775 ;
      LAYER CUT12 ;
        RECT 0.23 1.845 0.33 1.945 ;
        RECT 0.45 1.845 0.55 1.945 ;
        RECT 0.67 1.845 0.77 1.945 ;
        RECT 0.89 1.845 0.99 1.945 ;
        RECT 1.11 1.845 1.21 1.945 ;
        RECT 1.33 1.845 1.43 1.945 ;
        RECT 1.55 1.845 1.65 1.945 ;
        RECT 1.77 1.845 1.87 1.945 ;
        RECT 1.99 1.845 2.09 1.945 ;
        RECT 2.12 2.145 2.22 2.245 ;
        RECT 2.12 1.515 2.22 1.615 ;
        RECT 2.12 1.295 2.22 1.395 ;
        RECT 2.12 1.075 2.22 1.175 ;
        RECT 2.21 1.845 2.31 1.945 ;
        RECT 2.43 1.845 2.53 1.945 ;
        RECT 2.65 1.845 2.75 1.945 ;
        RECT 2.86 2.145 2.96 2.245 ;
        RECT 2.86 1.515 2.96 1.615 ;
        RECT 2.86 1.295 2.96 1.395 ;
        RECT 2.86 1.075 2.96 1.175 ;
        RECT 2.87 1.845 2.97 1.945 ;
        RECT 3.09 1.845 3.19 1.945 ;
        RECT 3.31 1.845 3.41 1.945 ;
        RECT 3.53 1.845 3.63 1.945 ;
        RECT 3.6 2.145 3.7 2.245 ;
        RECT 3.6 1.515 3.7 1.615 ;
        RECT 3.6 1.295 3.7 1.395 ;
        RECT 3.6 1.075 3.7 1.175 ;
        RECT 3.75 1.845 3.85 1.945 ;
        RECT 3.97 1.845 4.07 1.945 ;
        RECT 4.19 1.845 4.29 1.945 ;
        RECT 4.34 2.145 4.44 2.245 ;
        RECT 4.34 1.515 4.44 1.615 ;
        RECT 4.34 1.295 4.44 1.395 ;
        RECT 4.34 1.075 4.44 1.175 ;
        RECT 4.41 1.845 4.51 1.945 ;
        RECT 4.63 1.845 4.73 1.945 ;
        RECT 4.85 1.845 4.95 1.945 ;
        RECT 5.07 1.845 5.17 1.945 ;
        RECT 5.08 2.145 5.18 2.245 ;
        RECT 5.08 1.515 5.18 1.615 ;
        RECT 5.08 1.295 5.18 1.395 ;
        RECT 5.08 1.075 5.18 1.175 ;
        RECT 5.29 1.845 5.39 1.945 ;
        RECT 5.51 1.845 5.61 1.945 ;
        RECT 5.73 1.845 5.83 1.945 ;
        RECT 5.82 2.145 5.92 2.245 ;
        RECT 5.82 1.515 5.92 1.615 ;
        RECT 5.82 1.295 5.92 1.395 ;
        RECT 5.82 1.075 5.92 1.175 ;
        RECT 5.95 1.845 6.05 1.945 ;
        RECT 6.17 1.845 6.27 1.945 ;
        RECT 6.39 1.845 6.49 1.945 ;
        RECT 6.56 2.145 6.66 2.245 ;
        RECT 6.56 1.515 6.66 1.615 ;
        RECT 6.56 1.295 6.66 1.395 ;
        RECT 6.56 1.075 6.66 1.175 ;
        RECT 6.61 1.845 6.71 1.945 ;
        RECT 6.83 1.845 6.93 1.945 ;
        RECT 7.05 1.845 7.15 1.945 ;
        RECT 7.27 1.845 7.37 1.945 ;
        RECT 7.3 2.145 7.4 2.245 ;
        RECT 7.3 1.515 7.4 1.615 ;
        RECT 7.3 1.295 7.4 1.395 ;
    END
  END VDD
  PIN VDDSRC
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 0.08 2.41 9.72 3.01 ;
        RECT 0.08 0.31 9.72 0.91 ;
      LAYER CUT12 ;
        RECT 1.75 2.88 1.85 2.98 ;
        RECT 1.75 2.66 1.85 2.76 ;
        RECT 1.75 2.44 1.85 2.54 ;
        RECT 1.75 0.78 1.85 0.88 ;
        RECT 1.75 0.56 1.85 0.66 ;
        RECT 1.75 0.34 1.85 0.44 ;
        RECT 2.49 2.88 2.59 2.98 ;
        RECT 2.49 2.66 2.59 2.76 ;
        RECT 2.49 2.44 2.59 2.54 ;
        RECT 2.49 0.78 2.59 0.88 ;
        RECT 2.49 0.56 2.59 0.66 ;
        RECT 2.49 0.34 2.59 0.44 ;
        RECT 3.23 2.88 3.33 2.98 ;
        RECT 3.23 2.66 3.33 2.76 ;
        RECT 3.23 2.44 3.33 2.54 ;
        RECT 3.23 0.78 3.33 0.88 ;
        RECT 3.23 0.56 3.33 0.66 ;
        RECT 3.23 0.34 3.33 0.44 ;
        RECT 3.97 2.88 4.07 2.98 ;
        RECT 3.97 2.66 4.07 2.76 ;
        RECT 3.97 2.44 4.07 2.54 ;
        RECT 3.97 0.78 4.07 0.88 ;
        RECT 3.97 0.56 4.07 0.66 ;
        RECT 3.97 0.34 4.07 0.44 ;
        RECT 4.71 2.88 4.81 2.98 ;
        RECT 4.71 2.66 4.81 2.76 ;
        RECT 4.71 2.44 4.81 2.54 ;
        RECT 4.71 0.78 4.81 0.88 ;
        RECT 4.71 0.56 4.81 0.66 ;
        RECT 4.71 0.34 4.81 0.44 ;
        RECT 5.45 2.88 5.55 2.98 ;
        RECT 5.45 2.66 5.55 2.76 ;
        RECT 5.45 2.44 5.55 2.54 ;
        RECT 5.45 0.78 5.55 0.88 ;
        RECT 5.45 0.56 5.55 0.66 ;
        RECT 5.45 0.34 5.55 0.44 ;
        RECT 6.19 2.88 6.29 2.98 ;
        RECT 6.19 2.66 6.29 2.76 ;
        RECT 6.19 2.44 6.29 2.54 ;
        RECT 6.19 0.78 6.29 0.88 ;
        RECT 6.19 0.56 6.29 0.66 ;
        RECT 6.19 0.34 6.29 0.44 ;
        RECT 6.93 2.88 7.03 2.98 ;
        RECT 6.93 2.66 7.03 2.76 ;
        RECT 6.93 2.44 7.03 2.54 ;
        RECT 6.93 0.78 7.03 0.88 ;
        RECT 6.93 0.56 7.03 0.66 ;
        RECT 6.93 0.34 7.03 0.44 ;
        RECT 7.67 2.88 7.77 2.98 ;
        RECT 7.67 2.66 7.77 2.76 ;
        RECT 7.67 2.44 7.77 2.54 ;
        RECT 7.67 0.78 7.77 0.88 ;
        RECT 7.67 0.56 7.77 0.66 ;
        RECT 7.67 0.34 7.77 0.44 ;
        RECT 7.95 2.88 8.05 2.98 ;
        RECT 7.95 2.66 8.05 2.76 ;
        RECT 7.95 2.44 8.05 2.54 ;
        RECT 7.95 0.78 8.05 0.88 ;
        RECT 7.95 0.56 8.05 0.66 ;
        RECT 7.95 0.34 8.05 0.44 ;
    END
  END VDDSRC
  OBS
    LAYER MET1 ;
      RECT 1.73 2.08 1.87 3.07 ;
      RECT 1.73 0.28 1.87 1.52 ;
      RECT 2.1 1.96 2.24 3.07 ;
      RECT 2.1 0.28 2.24 1.64 ;
      RECT 2.47 2.08 2.61 3.07 ;
      RECT 2.47 0.28 2.61 1.52 ;
      RECT 2.84 1.96 2.98 3.07 ;
      RECT 2.84 0.28 2.98 1.64 ;
      RECT 3.21 2.08 3.35 3.07 ;
      RECT 3.21 0.28 3.35 1.52 ;
      RECT 3.58 1.96 3.72 3.07 ;
      RECT 3.58 0.28 3.72 1.64 ;
      RECT 3.95 2.08 4.09 3.07 ;
      RECT 3.95 0.28 4.09 1.52 ;
      RECT 4.32 1.96 4.46 3.07 ;
      RECT 4.32 0.28 4.46 1.64 ;
      RECT 4.69 2.08 4.83 3.07 ;
      RECT 4.69 0.28 4.83 1.52 ;
      RECT 5.06 1.96 5.2 3.07 ;
      RECT 5.06 0.28 5.2 1.64 ;
      RECT 5.43 2.08 5.57 3.07 ;
      RECT 5.43 0.28 5.57 1.52 ;
      RECT 5.8 1.96 5.94 3.07 ;
      RECT 5.8 0.28 5.94 1.64 ;
      RECT 6.17 2.08 6.31 3.07 ;
      RECT 6.17 0.28 6.31 1.52 ;
      RECT 6.54 1.96 6.68 3.07 ;
      RECT 6.54 0.28 6.68 1.64 ;
      RECT 6.91 2.08 7.05 3.07 ;
      RECT 6.91 0.28 7.05 1.52 ;
      RECT 7.28 1.96 7.42 3.07 ;
      RECT 7.28 0.28 7.42 1.64 ;
      RECT 7.65 2.08 7.79 3.07 ;
      RECT 7.65 0.28 7.79 1.52 ;
      RECT 7.93 2.08 8.07 3.07 ;
      RECT 7.93 0.28 8.07 1.52 ;
  END
END DSIPGX2LPSCCS1

MACRO DSIPGX2LCNRC1
  CLASS RING ;
  ORIGIN 0 0 ;
  FOREIGN DSIPGX2LCNRC1 0 0 ;
  SIZE 11.57 BY 11.57 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0.23 0.23 0.37 11.57 ;
        RECT 0.23 0.23 11.57 0.37 ;
      LAYER CUT01 ;
        RECT 0.255 11.255 0.345 11.345 ;
        RECT 0.255 11.035 0.345 11.125 ;
        RECT 0.255 10.815 0.345 10.905 ;
        RECT 0.255 10.595 0.345 10.685 ;
        RECT 0.255 10.375 0.345 10.465 ;
        RECT 0.255 10.155 0.345 10.245 ;
        RECT 0.255 9.935 0.345 10.025 ;
        RECT 0.255 9.715 0.345 9.805 ;
        RECT 0.255 9.495 0.345 9.585 ;
        RECT 0.255 9.275 0.345 9.365 ;
        RECT 0.255 9.055 0.345 9.145 ;
        RECT 0.255 8.835 0.345 8.925 ;
        RECT 0.255 8.615 0.345 8.705 ;
        RECT 0.255 8.395 0.345 8.485 ;
        RECT 0.255 8.175 0.345 8.265 ;
        RECT 0.255 7.955 0.345 8.045 ;
        RECT 0.255 7.735 0.345 7.825 ;
        RECT 0.255 7.515 0.345 7.605 ;
        RECT 0.255 7.295 0.345 7.385 ;
        RECT 0.255 7.075 0.345 7.165 ;
        RECT 0.255 6.855 0.345 6.945 ;
        RECT 0.255 6.635 0.345 6.725 ;
        RECT 0.255 6.415 0.345 6.505 ;
        RECT 0.255 6.195 0.345 6.285 ;
        RECT 0.255 5.975 0.345 6.065 ;
        RECT 0.255 5.755 0.345 5.845 ;
        RECT 0.255 5.535 0.345 5.625 ;
        RECT 0.255 5.315 0.345 5.405 ;
        RECT 0.255 5.095 0.345 5.185 ;
        RECT 0.255 4.875 0.345 4.965 ;
        RECT 0.255 4.655 0.345 4.745 ;
        RECT 0.255 4.435 0.345 4.525 ;
        RECT 0.255 4.215 0.345 4.305 ;
        RECT 0.255 3.995 0.345 4.085 ;
        RECT 0.255 3.775 0.345 3.865 ;
        RECT 0.255 3.555 0.345 3.645 ;
        RECT 0.255 3.335 0.345 3.425 ;
        RECT 0.255 3.115 0.345 3.205 ;
        RECT 0.255 2.895 0.345 2.985 ;
        RECT 0.255 2.675 0.345 2.765 ;
        RECT 0.255 2.455 0.345 2.545 ;
        RECT 0.255 2.235 0.345 2.325 ;
        RECT 0.255 2.015 0.345 2.105 ;
        RECT 0.255 1.795 0.345 1.885 ;
        RECT 0.255 1.575 0.345 1.665 ;
        RECT 0.255 1.355 0.345 1.445 ;
        RECT 0.255 1.135 0.345 1.225 ;
        RECT 0.255 0.915 0.345 1.005 ;
        RECT 0.255 0.695 0.345 0.785 ;
        RECT 0.255 0.475 0.345 0.565 ;
        RECT 0.475 0.255 0.565 0.345 ;
        RECT 0.695 0.255 0.785 0.345 ;
        RECT 0.915 0.255 1.005 0.345 ;
        RECT 1.135 0.255 1.225 0.345 ;
        RECT 1.355 0.255 1.445 0.345 ;
        RECT 1.575 0.255 1.665 0.345 ;
        RECT 1.795 0.255 1.885 0.345 ;
        RECT 2.015 0.255 2.105 0.345 ;
        RECT 2.235 0.255 2.325 0.345 ;
        RECT 2.455 0.255 2.545 0.345 ;
        RECT 2.675 0.255 2.765 0.345 ;
        RECT 2.895 0.255 2.985 0.345 ;
        RECT 3.115 0.255 3.205 0.345 ;
        RECT 3.335 0.255 3.425 0.345 ;
        RECT 3.555 0.255 3.645 0.345 ;
        RECT 3.775 0.255 3.865 0.345 ;
        RECT 3.995 0.255 4.085 0.345 ;
        RECT 4.215 0.255 4.305 0.345 ;
        RECT 4.435 0.255 4.525 0.345 ;
        RECT 4.655 0.255 4.745 0.345 ;
        RECT 4.875 0.255 4.965 0.345 ;
        RECT 5.095 0.255 5.185 0.345 ;
        RECT 5.315 0.255 5.405 0.345 ;
        RECT 5.535 0.255 5.625 0.345 ;
        RECT 5.755 0.255 5.845 0.345 ;
        RECT 5.975 0.255 6.065 0.345 ;
        RECT 6.195 0.255 6.285 0.345 ;
        RECT 6.415 0.255 6.505 0.345 ;
        RECT 6.635 0.255 6.725 0.345 ;
        RECT 6.855 0.255 6.945 0.345 ;
        RECT 7.075 0.255 7.165 0.345 ;
        RECT 7.295 0.255 7.385 0.345 ;
        RECT 7.515 0.255 7.605 0.345 ;
        RECT 7.735 0.255 7.825 0.345 ;
        RECT 7.955 0.255 8.045 0.345 ;
        RECT 8.175 0.255 8.265 0.345 ;
        RECT 8.395 0.255 8.485 0.345 ;
        RECT 8.615 0.255 8.705 0.345 ;
        RECT 8.835 0.255 8.925 0.345 ;
        RECT 9.055 0.255 9.145 0.345 ;
        RECT 9.275 0.255 9.365 0.345 ;
        RECT 9.495 0.255 9.585 0.345 ;
        RECT 9.715 0.255 9.805 0.345 ;
        RECT 9.935 0.255 10.025 0.345 ;
        RECT 10.155 0.255 10.245 0.345 ;
        RECT 10.375 0.255 10.465 0.345 ;
        RECT 10.595 0.255 10.685 0.345 ;
        RECT 10.815 0.255 10.905 0.345 ;
        RECT 11.035 0.255 11.125 0.345 ;
        RECT 11.255 0.255 11.345 0.345 ;
    END
  END VSS
  PIN VDDPD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 9.81 9.81 11.25 11.57 ;
        RECT 9.81 9.81 11.57 11.25 ;
        RECT 8.22 8.22 9.66 11.57 ;
        RECT 8.22 8.22 11.57 9.66 ;
        RECT 6.63 6.63 8.07 11.57 ;
        RECT 6.63 6.63 11.57 8.07 ;
    END
  END VDDPD
  PIN VDDSRC
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 3.79 3.79 11.57 5.23 ;
        RECT 2.2 2.2 3.64 11.57 ;
        RECT 2.2 2.2 11.57 3.64 ;
        RECT 0.61 0.61 2.05 11.57 ;
        RECT 0.61 0.61 11.57 2.05 ;
      LAYER CUT12 ;
        RECT 1.28 1.28 1.38 1.38 ;
        RECT 1.5 1.28 1.6 1.38 ;
        RECT 1.72 1.28 1.82 1.38 ;
        RECT 1.94 1.28 2.04 1.38 ;
      LAYER CUT01 ;
        RECT 1.285 1.285 1.375 1.375 ;
        RECT 1.505 1.285 1.595 1.375 ;
        RECT 1.725 1.285 1.815 1.375 ;
        RECT 1.945 1.285 2.035 1.375 ;
      LAYER MET1 ;
        RECT 1.235 1.26 2.085 1.4 ;
      LAYER MET2 ;
        RECT 3.79 3.79 5.23 11.57 ;
    END
  END VDDSRC
END DSIPGX2LCNRC1
MACRO DSIPGX2LCNRC2
  CLASS RING ;
  ORIGIN 0 0 ;
  FOREIGN DSIPGX2LCNRC2 0 0 ;
  SIZE 11.57 BY 11.57 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 11.2 11.2 11.34 11.57 ;
        RECT 11.2 11.2 11.57 11.34 ;
      LAYER CUT01 ;
        RECT 11.25 11.225 11.34 11.315 ;
    END
  END VSS
  PIN VDDPD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 3.5 3.5 4.94 11.57 ;
        RECT 3.5 3.5 11.57 4.94 ;
        RECT 1.91 1.91 3.35 11.57 ;
        RECT 1.91 1.91 11.57 3.35 ;
        RECT 0.32 0.32 1.76 11.57 ;
        RECT 0.32 0.32 11.57 1.76 ;
    END
  END VDDPD
  PIN VDDSRC
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 10.145 10.17 10.995 10.31 ;
      LAYER MET2 ;
        RECT 9.52 9.52 10.96 11.57 ;
        RECT 9.52 9.52 11.57 10.96 ;
        RECT 7.93 7.93 9.37 11.57 ;
        RECT 7.93 7.93 11.57 9.37 ;
        RECT 6.34 6.34 7.78 11.57 ;
        RECT 6.34 6.34 11.57 7.78 ;
      LAYER CUT12 ;
        RECT 10.19 10.19 10.29 10.29 ;
        RECT 10.41 10.19 10.51 10.29 ;
        RECT 10.63 10.19 10.73 10.29 ;
        RECT 10.85 10.19 10.95 10.29 ;
      LAYER CUT01 ;
        RECT 10.195 10.195 10.285 10.285 ;
        RECT 10.415 10.195 10.505 10.285 ;
        RECT 10.635 10.195 10.725 10.285 ;
        RECT 10.855 10.195 10.945 10.285 ;
    END
  END VDDSRC
END DSIPGX2LCNRC2
MACRO DSIPGX2LPSRCL1
  CLASS RING ;
  ORIGIN 0 0 ;
  FOREIGN DSIPGX2LPSRCL1 0 0 ;
  SIZE 7.68 BY 11.57 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 0.23 7.68 0.37 ;
      LAYER CUT01 ;
        RECT 0.52 0.255 0.61 0.345 ;
        RECT 0.74 0.255 0.83 0.345 ;
        RECT 0.96 0.255 1.05 0.345 ;
        RECT 1.18 0.255 1.27 0.345 ;
        RECT 1.4 0.255 1.49 0.345 ;
        RECT 1.62 0.255 1.71 0.345 ;
        RECT 1.84 0.255 1.93 0.345 ;
        RECT 2.06 0.255 2.15 0.345 ;
        RECT 2.28 0.255 2.37 0.345 ;
        RECT 2.5 0.255 2.59 0.345 ;
        RECT 2.72 0.255 2.81 0.345 ;
        RECT 2.94 0.255 3.03 0.345 ;
        RECT 3.16 0.255 3.25 0.345 ;
        RECT 3.38 0.255 3.47 0.345 ;
        RECT 3.6 0.255 3.69 0.345 ;
        RECT 3.82 0.255 3.91 0.345 ;
        RECT 4.04 0.255 4.13 0.345 ;
        RECT 4.26 0.255 4.35 0.345 ;
        RECT 4.48 0.255 4.57 0.345 ;
        RECT 4.7 0.255 4.79 0.345 ;
        RECT 4.92 0.255 5.01 0.345 ;
        RECT 5.14 0.255 5.23 0.345 ;
        RECT 5.36 0.255 5.45 0.345 ;
        RECT 5.58 0.255 5.67 0.345 ;
        RECT 5.8 0.255 5.89 0.345 ;
        RECT 6.02 0.255 6.11 0.345 ;
        RECT 6.24 0.255 6.33 0.345 ;
        RECT 6.46 0.255 6.55 0.345 ;
        RECT 6.68 0.255 6.77 0.345 ;
        RECT 6.9 0.255 6.99 0.345 ;
        RECT 7.12 0.255 7.21 0.345 ;
        RECT 7.34 0.255 7.43 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE ANALOG ;
      ANTENNAGATEAREA 30.4 LAYER MET1 ;
      ANTENNAGATEAREA 30.4 LAYER MET2 ;
    ANTENNAMAXCUTCAR 3.552632 LAYER CUT01 ;
    SUPPLYSENSITIVITY VDDSRC ;
    GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 0.15 5.38 0.29 11.16 ;
        RECT 0.15 11.02 7.36 11.16 ;
      LAYER MET2 ;
        RECT 0.15 5.38 0.29 6.48 ;
      LAYER CUT12 ;
        RECT 0.17 6.34 0.27 6.44 ;
        RECT 0.17 6.11 0.27 6.21 ;
        RECT 0.17 5.88 0.27 5.98 ;
        RECT 0.17 5.65 0.27 5.75 ;
        RECT 0.17 5.42 0.27 5.52 ;
      LAYER CUT01 ;
        RECT 0.63 11.045 0.72 11.135 ;
        RECT 0.85 11.045 0.94 11.135 ;
        RECT 1.07 11.045 1.16 11.135 ;
        RECT 1.29 11.045 1.38 11.135 ;
        RECT 1.51 11.045 1.6 11.135 ;
        RECT 1.73 11.045 1.82 11.135 ;
        RECT 1.95 11.045 2.04 11.135 ;
        RECT 2.17 11.045 2.26 11.135 ;
        RECT 2.39 11.045 2.48 11.135 ;
        RECT 2.61 11.045 2.7 11.135 ;
        RECT 2.83 11.045 2.92 11.135 ;
        RECT 3.05 11.045 3.14 11.135 ;
        RECT 3.27 11.045 3.36 11.135 ;
        RECT 3.49 11.045 3.58 11.135 ;
        RECT 3.71 11.045 3.8 11.135 ;
        RECT 3.93 11.045 4.02 11.135 ;
        RECT 4.15 11.045 4.24 11.135 ;
        RECT 4.37 11.045 4.46 11.135 ;
        RECT 4.59 11.045 4.68 11.135 ;
        RECT 4.81 11.045 4.9 11.135 ;
        RECT 5.03 11.045 5.12 11.135 ;
        RECT 5.25 11.045 5.34 11.135 ;
        RECT 5.47 11.045 5.56 11.135 ;
        RECT 5.69 11.045 5.78 11.135 ;
        RECT 5.91 11.045 6 11.135 ;
        RECT 6.13 11.045 6.22 11.135 ;
        RECT 6.35 11.045 6.44 11.135 ;
        RECT 6.57 11.045 6.66 11.135 ;
        RECT 6.79 11.045 6.88 11.135 ;
        RECT 7.01 11.045 7.1 11.135 ;
        RECT 7.23 11.045 7.32 11.135 ;
    END
  END A
  PIN VDDPD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER CUT12 ;
        RECT 6.7 8.545 6.8 8.645 ;
        RECT 6.7 8.315 6.8 8.415 ;
        RECT 6.7 7.875 6.8 7.975 ;
        RECT 6.7 7.645 6.8 7.745 ;
        RECT 6.7 7.415 6.8 7.515 ;
        RECT 6.7 7.185 6.8 7.285 ;
        RECT 6.7 6.955 6.8 7.055 ;
        RECT 6.7 6.725 6.8 6.825 ;
        RECT 7.44 10.765 7.54 10.865 ;
        RECT 7.44 10.535 7.54 10.635 ;
        RECT 7.44 10.305 7.54 10.405 ;
        RECT 7.44 10.075 7.54 10.175 ;
        RECT 7.44 9.845 7.54 9.945 ;
        RECT 7.44 9.465 7.54 9.565 ;
        RECT 7.44 9.235 7.54 9.335 ;
        RECT 7.44 9.005 7.54 9.105 ;
        RECT 7.44 8.775 7.54 8.875 ;
        RECT 7.44 8.545 7.54 8.645 ;
        RECT 7.44 8.315 7.54 8.415 ;
        RECT 7.44 7.875 7.54 7.975 ;
        RECT 7.44 7.645 7.54 7.745 ;
        RECT 7.44 7.415 7.54 7.515 ;
        RECT 7.44 7.185 7.54 7.285 ;
        RECT 7.44 6.955 7.54 7.055 ;
        RECT 7.44 6.725 7.54 6.825 ;
      LAYER MET2 ;
        RECT 0 9.81 7.68 11.25 ;
        RECT 0 8.22 7.68 9.66 ;
        RECT 0 6.63 7.68 8.07 ;
      LAYER CUT12 ;
        RECT 0.78 10.765 0.88 10.865 ;
        RECT 0.78 10.535 0.88 10.635 ;
        RECT 0.78 10.305 0.88 10.405 ;
        RECT 0.78 10.075 0.88 10.175 ;
        RECT 0.78 9.845 0.88 9.945 ;
        RECT 0.78 9.465 0.88 9.565 ;
        RECT 0.78 9.235 0.88 9.335 ;
        RECT 0.78 9.005 0.88 9.105 ;
        RECT 0.78 8.775 0.88 8.875 ;
        RECT 0.78 8.545 0.88 8.645 ;
        RECT 0.78 8.315 0.88 8.415 ;
        RECT 0.78 7.875 0.88 7.975 ;
        RECT 0.78 7.645 0.88 7.745 ;
        RECT 0.78 7.415 0.88 7.515 ;
        RECT 0.78 7.185 0.88 7.285 ;
        RECT 0.78 6.955 0.88 7.055 ;
        RECT 0.78 6.725 0.88 6.825 ;
        RECT 1.52 10.765 1.62 10.865 ;
        RECT 1.52 10.535 1.62 10.635 ;
        RECT 1.52 10.305 1.62 10.405 ;
        RECT 1.52 10.075 1.62 10.175 ;
        RECT 1.52 9.845 1.62 9.945 ;
        RECT 1.52 9.465 1.62 9.565 ;
        RECT 1.52 9.235 1.62 9.335 ;
        RECT 1.52 9.005 1.62 9.105 ;
        RECT 1.52 8.775 1.62 8.875 ;
        RECT 1.52 8.545 1.62 8.645 ;
        RECT 1.52 8.315 1.62 8.415 ;
        RECT 1.52 7.875 1.62 7.975 ;
        RECT 1.52 7.645 1.62 7.745 ;
        RECT 1.52 7.415 1.62 7.515 ;
        RECT 1.52 7.185 1.62 7.285 ;
        RECT 1.52 6.955 1.62 7.055 ;
        RECT 1.52 6.725 1.62 6.825 ;
        RECT 2.26 10.765 2.36 10.865 ;
        RECT 2.26 10.535 2.36 10.635 ;
        RECT 2.26 10.305 2.36 10.405 ;
        RECT 2.26 10.075 2.36 10.175 ;
        RECT 2.26 9.845 2.36 9.945 ;
        RECT 2.26 9.465 2.36 9.565 ;
        RECT 2.26 9.235 2.36 9.335 ;
        RECT 2.26 9.005 2.36 9.105 ;
        RECT 2.26 8.775 2.36 8.875 ;
        RECT 2.26 8.545 2.36 8.645 ;
        RECT 2.26 8.315 2.36 8.415 ;
        RECT 2.26 7.875 2.36 7.975 ;
        RECT 2.26 7.645 2.36 7.745 ;
        RECT 2.26 7.415 2.36 7.515 ;
        RECT 2.26 7.185 2.36 7.285 ;
        RECT 2.26 6.955 2.36 7.055 ;
        RECT 2.26 6.725 2.36 6.825 ;
        RECT 3 10.765 3.1 10.865 ;
        RECT 3 10.535 3.1 10.635 ;
        RECT 3 10.305 3.1 10.405 ;
        RECT 3 10.075 3.1 10.175 ;
        RECT 3 9.845 3.1 9.945 ;
        RECT 3 9.465 3.1 9.565 ;
        RECT 3 9.235 3.1 9.335 ;
        RECT 3 9.005 3.1 9.105 ;
        RECT 3 8.775 3.1 8.875 ;
        RECT 3 8.545 3.1 8.645 ;
        RECT 3 8.315 3.1 8.415 ;
        RECT 3 7.875 3.1 7.975 ;
        RECT 3 7.645 3.1 7.745 ;
        RECT 3 7.415 3.1 7.515 ;
        RECT 3 7.185 3.1 7.285 ;
        RECT 3 6.955 3.1 7.055 ;
        RECT 3 6.725 3.1 6.825 ;
        RECT 3.74 10.765 3.84 10.865 ;
        RECT 3.74 10.535 3.84 10.635 ;
        RECT 3.74 10.305 3.84 10.405 ;
        RECT 3.74 10.075 3.84 10.175 ;
        RECT 3.74 9.845 3.84 9.945 ;
        RECT 3.74 9.465 3.84 9.565 ;
        RECT 3.74 9.235 3.84 9.335 ;
        RECT 3.74 9.005 3.84 9.105 ;
        RECT 3.74 8.775 3.84 8.875 ;
        RECT 3.74 8.545 3.84 8.645 ;
        RECT 3.74 8.315 3.84 8.415 ;
        RECT 3.74 7.875 3.84 7.975 ;
        RECT 3.74 7.645 3.84 7.745 ;
        RECT 3.74 7.415 3.84 7.515 ;
        RECT 3.74 7.185 3.84 7.285 ;
        RECT 3.74 6.955 3.84 7.055 ;
        RECT 3.74 6.725 3.84 6.825 ;
        RECT 4.48 10.765 4.58 10.865 ;
        RECT 4.48 10.535 4.58 10.635 ;
        RECT 4.48 10.305 4.58 10.405 ;
        RECT 4.48 10.075 4.58 10.175 ;
        RECT 4.48 9.845 4.58 9.945 ;
        RECT 4.48 9.465 4.58 9.565 ;
        RECT 4.48 9.235 4.58 9.335 ;
        RECT 4.48 9.005 4.58 9.105 ;
        RECT 4.48 8.775 4.58 8.875 ;
        RECT 4.48 8.545 4.58 8.645 ;
        RECT 4.48 8.315 4.58 8.415 ;
        RECT 4.48 7.875 4.58 7.975 ;
        RECT 4.48 7.645 4.58 7.745 ;
        RECT 4.48 7.415 4.58 7.515 ;
        RECT 4.48 7.185 4.58 7.285 ;
        RECT 4.48 6.955 4.58 7.055 ;
        RECT 4.48 6.725 4.58 6.825 ;
        RECT 5.22 10.765 5.32 10.865 ;
        RECT 5.22 10.535 5.32 10.635 ;
        RECT 5.22 10.305 5.32 10.405 ;
        RECT 5.22 10.075 5.32 10.175 ;
        RECT 5.22 9.845 5.32 9.945 ;
        RECT 5.22 9.465 5.32 9.565 ;
        RECT 5.22 9.235 5.32 9.335 ;
        RECT 5.22 9.005 5.32 9.105 ;
        RECT 5.22 8.775 5.32 8.875 ;
        RECT 5.22 8.545 5.32 8.645 ;
        RECT 5.22 8.315 5.32 8.415 ;
        RECT 5.22 7.875 5.32 7.975 ;
        RECT 5.22 7.645 5.32 7.745 ;
        RECT 5.22 7.415 5.32 7.515 ;
        RECT 5.22 7.185 5.32 7.285 ;
        RECT 5.22 6.955 5.32 7.055 ;
        RECT 5.22 6.725 5.32 6.825 ;
        RECT 5.96 10.765 6.06 10.865 ;
        RECT 5.96 10.535 6.06 10.635 ;
        RECT 5.96 10.305 6.06 10.405 ;
        RECT 5.96 10.075 6.06 10.175 ;
        RECT 5.96 9.845 6.06 9.945 ;
        RECT 5.96 9.465 6.06 9.565 ;
        RECT 5.96 9.235 6.06 9.335 ;
        RECT 5.96 9.005 6.06 9.105 ;
        RECT 5.96 8.775 6.06 8.875 ;
        RECT 5.96 8.545 6.06 8.645 ;
        RECT 5.96 8.315 6.06 8.415 ;
        RECT 5.96 7.875 6.06 7.975 ;
        RECT 5.96 7.645 6.06 7.745 ;
        RECT 5.96 7.415 6.06 7.515 ;
        RECT 5.96 7.185 6.06 7.285 ;
        RECT 5.96 6.955 6.06 7.055 ;
        RECT 5.96 6.725 6.06 6.825 ;
        RECT 6.7 10.765 6.8 10.865 ;
        RECT 6.7 10.535 6.8 10.635 ;
        RECT 6.7 10.305 6.8 10.405 ;
        RECT 6.7 10.075 6.8 10.175 ;
        RECT 6.7 9.845 6.8 9.945 ;
        RECT 6.7 9.465 6.8 9.565 ;
        RECT 6.7 9.235 6.8 9.335 ;
        RECT 6.7 9.005 6.8 9.105 ;
        RECT 6.7 8.775 6.8 8.875 ;
    END
  END VDDPD
  PIN VDDSRC
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 0 3.79 7.68 5.23 ;
        RECT 0 2.2 7.68 3.64 ;
        RECT 0 0.61 7.68 2.05 ;
      LAYER CUT12 ;
        RECT 0.41 5.035 0.51 5.135 ;
        RECT 0.41 4.805 0.51 4.905 ;
        RECT 0.41 4.575 0.51 4.675 ;
        RECT 0.41 4.345 0.51 4.445 ;
        RECT 0.41 4.115 0.51 4.215 ;
        RECT 0.41 3.885 0.51 3.985 ;
        RECT 0.41 3.445 0.51 3.545 ;
        RECT 0.41 3.215 0.51 3.315 ;
        RECT 0.41 2.985 0.51 3.085 ;
        RECT 0.41 2.755 0.51 2.855 ;
        RECT 0.41 2.525 0.51 2.625 ;
        RECT 0.41 2.295 0.51 2.395 ;
        RECT 0.41 1.855 0.51 1.955 ;
        RECT 0.41 1.625 0.51 1.725 ;
        RECT 0.41 1.395 0.51 1.495 ;
        RECT 0.41 1.165 0.51 1.265 ;
        RECT 0.41 0.935 0.51 1.035 ;
        RECT 0.48 0.65 0.58 0.75 ;
        RECT 0.71 0.65 0.81 0.75 ;
        RECT 0.94 0.65 1.04 0.75 ;
        RECT 1.15 5.035 1.25 5.135 ;
        RECT 1.15 4.805 1.25 4.905 ;
        RECT 1.15 4.575 1.25 4.675 ;
        RECT 1.15 4.345 1.25 4.445 ;
        RECT 1.15 4.115 1.25 4.215 ;
        RECT 1.15 3.885 1.25 3.985 ;
        RECT 1.15 3.445 1.25 3.545 ;
        RECT 1.15 3.215 1.25 3.315 ;
        RECT 1.15 2.985 1.25 3.085 ;
        RECT 1.15 2.755 1.25 2.855 ;
        RECT 1.15 2.525 1.25 2.625 ;
        RECT 1.15 2.295 1.25 2.395 ;
        RECT 1.15 1.855 1.25 1.955 ;
        RECT 1.15 1.625 1.25 1.725 ;
        RECT 1.15 1.395 1.25 1.495 ;
        RECT 1.15 1.165 1.25 1.265 ;
        RECT 1.15 0.935 1.25 1.035 ;
        RECT 1.17 0.65 1.27 0.75 ;
        RECT 1.4 0.65 1.5 0.75 ;
        RECT 1.63 0.65 1.73 0.75 ;
        RECT 1.86 0.65 1.96 0.75 ;
        RECT 1.89 5.035 1.99 5.135 ;
        RECT 1.89 4.805 1.99 4.905 ;
        RECT 1.89 4.575 1.99 4.675 ;
        RECT 1.89 4.345 1.99 4.445 ;
        RECT 1.89 4.115 1.99 4.215 ;
        RECT 1.89 3.885 1.99 3.985 ;
        RECT 1.89 3.445 1.99 3.545 ;
        RECT 1.89 3.215 1.99 3.315 ;
        RECT 1.89 2.985 1.99 3.085 ;
        RECT 1.89 2.755 1.99 2.855 ;
        RECT 1.89 2.525 1.99 2.625 ;
        RECT 1.89 2.295 1.99 2.395 ;
        RECT 1.89 1.855 1.99 1.955 ;
        RECT 1.89 1.625 1.99 1.725 ;
        RECT 1.89 1.395 1.99 1.495 ;
        RECT 1.89 1.165 1.99 1.265 ;
        RECT 1.89 0.935 1.99 1.035 ;
        RECT 2.09 0.65 2.19 0.75 ;
        RECT 2.32 0.65 2.42 0.75 ;
        RECT 2.55 0.65 2.65 0.75 ;
        RECT 2.63 5.035 2.73 5.135 ;
        RECT 2.63 4.805 2.73 4.905 ;
        RECT 2.63 4.575 2.73 4.675 ;
        RECT 2.63 4.345 2.73 4.445 ;
        RECT 2.63 4.115 2.73 4.215 ;
        RECT 2.63 3.885 2.73 3.985 ;
        RECT 2.63 3.445 2.73 3.545 ;
        RECT 2.63 3.215 2.73 3.315 ;
        RECT 2.63 2.985 2.73 3.085 ;
        RECT 2.63 2.755 2.73 2.855 ;
        RECT 2.63 2.525 2.73 2.625 ;
        RECT 2.63 2.295 2.73 2.395 ;
        RECT 2.63 1.855 2.73 1.955 ;
        RECT 2.63 1.625 2.73 1.725 ;
        RECT 2.63 1.395 2.73 1.495 ;
        RECT 2.63 1.165 2.73 1.265 ;
        RECT 2.63 0.935 2.73 1.035 ;
        RECT 2.78 0.65 2.88 0.75 ;
        RECT 3.01 0.65 3.11 0.75 ;
        RECT 3.24 0.65 3.34 0.75 ;
        RECT 3.37 5.035 3.47 5.135 ;
        RECT 7.07 2.525 7.17 2.625 ;
        RECT 7.07 2.295 7.17 2.395 ;
        RECT 7.07 1.855 7.17 1.955 ;
        RECT 7.07 1.625 7.17 1.725 ;
        RECT 7.07 1.395 7.17 1.495 ;
        RECT 7.07 1.165 7.17 1.265 ;
        RECT 7.07 0.935 7.17 1.035 ;
        RECT 7.15 0.65 7.25 0.75 ;
        RECT 7.38 0.65 7.48 0.75 ;
        RECT 3.37 4.805 3.47 4.905 ;
        RECT 3.37 4.575 3.47 4.675 ;
        RECT 3.37 4.345 3.47 4.445 ;
        RECT 3.37 4.115 3.47 4.215 ;
        RECT 3.37 3.885 3.47 3.985 ;
        RECT 3.37 3.445 3.47 3.545 ;
        RECT 3.37 3.215 3.47 3.315 ;
        RECT 3.37 2.985 3.47 3.085 ;
        RECT 3.37 2.755 3.47 2.855 ;
        RECT 3.37 2.525 3.47 2.625 ;
        RECT 3.37 2.295 3.47 2.395 ;
        RECT 3.37 1.855 3.47 1.955 ;
        RECT 3.37 1.625 3.47 1.725 ;
        RECT 3.37 1.395 3.47 1.495 ;
        RECT 3.37 1.165 3.47 1.265 ;
        RECT 3.37 0.935 3.47 1.035 ;
        RECT 3.47 0.65 3.57 0.75 ;
        RECT 3.7 0.65 3.8 0.75 ;
        RECT 3.93 0.65 4.03 0.75 ;
        RECT 4.11 5.035 4.21 5.135 ;
        RECT 4.11 4.805 4.21 4.905 ;
        RECT 4.11 4.575 4.21 4.675 ;
        RECT 4.11 4.345 4.21 4.445 ;
        RECT 4.11 4.115 4.21 4.215 ;
        RECT 4.11 3.885 4.21 3.985 ;
        RECT 4.11 3.445 4.21 3.545 ;
        RECT 4.11 3.215 4.21 3.315 ;
        RECT 4.11 2.985 4.21 3.085 ;
        RECT 4.11 2.755 4.21 2.855 ;
        RECT 4.11 2.525 4.21 2.625 ;
        RECT 4.11 2.295 4.21 2.395 ;
        RECT 4.11 1.855 4.21 1.955 ;
        RECT 4.11 1.625 4.21 1.725 ;
        RECT 4.11 1.395 4.21 1.495 ;
        RECT 4.11 1.165 4.21 1.265 ;
        RECT 4.11 0.935 4.21 1.035 ;
        RECT 4.16 0.65 4.26 0.75 ;
        RECT 4.39 0.65 4.49 0.75 ;
        RECT 4.62 0.65 4.72 0.75 ;
        RECT 4.85 5.035 4.95 5.135 ;
        RECT 4.85 4.805 4.95 4.905 ;
        RECT 4.85 4.575 4.95 4.675 ;
        RECT 4.85 4.345 4.95 4.445 ;
        RECT 4.85 4.115 4.95 4.215 ;
        RECT 4.85 3.885 4.95 3.985 ;
        RECT 4.85 3.445 4.95 3.545 ;
        RECT 4.85 3.215 4.95 3.315 ;
        RECT 4.85 2.985 4.95 3.085 ;
        RECT 4.85 2.755 4.95 2.855 ;
        RECT 4.85 2.525 4.95 2.625 ;
        RECT 4.85 2.295 4.95 2.395 ;
        RECT 4.85 1.855 4.95 1.955 ;
        RECT 4.85 1.625 4.95 1.725 ;
        RECT 4.85 1.395 4.95 1.495 ;
        RECT 4.85 1.165 4.95 1.265 ;
        RECT 4.85 0.935 4.95 1.035 ;
        RECT 4.85 0.65 4.95 0.75 ;
        RECT 5.08 0.65 5.18 0.75 ;
        RECT 5.31 0.65 5.41 0.75 ;
        RECT 5.54 0.65 5.64 0.75 ;
        RECT 5.59 5.035 5.69 5.135 ;
        RECT 5.59 4.805 5.69 4.905 ;
        RECT 5.59 4.575 5.69 4.675 ;
        RECT 5.59 4.345 5.69 4.445 ;
        RECT 5.59 4.115 5.69 4.215 ;
        RECT 5.59 3.885 5.69 3.985 ;
        RECT 5.59 3.445 5.69 3.545 ;
        RECT 5.59 3.215 5.69 3.315 ;
        RECT 5.59 2.985 5.69 3.085 ;
        RECT 5.59 2.755 5.69 2.855 ;
        RECT 5.59 2.525 5.69 2.625 ;
        RECT 5.59 2.295 5.69 2.395 ;
        RECT 5.59 1.855 5.69 1.955 ;
        RECT 5.59 1.625 5.69 1.725 ;
        RECT 5.59 1.395 5.69 1.495 ;
        RECT 5.59 1.165 5.69 1.265 ;
        RECT 5.59 0.935 5.69 1.035 ;
        RECT 5.77 0.65 5.87 0.75 ;
        RECT 6 0.65 6.1 0.75 ;
        RECT 6.23 0.65 6.33 0.75 ;
        RECT 6.33 5.035 6.43 5.135 ;
        RECT 6.33 4.805 6.43 4.905 ;
        RECT 6.33 4.575 6.43 4.675 ;
        RECT 6.33 4.345 6.43 4.445 ;
        RECT 6.33 4.115 6.43 4.215 ;
        RECT 6.33 3.885 6.43 3.985 ;
        RECT 6.33 3.445 6.43 3.545 ;
        RECT 6.33 3.215 6.43 3.315 ;
        RECT 6.33 2.985 6.43 3.085 ;
        RECT 6.33 2.755 6.43 2.855 ;
        RECT 6.33 2.525 6.43 2.625 ;
        RECT 6.33 2.295 6.43 2.395 ;
        RECT 6.33 1.855 6.43 1.955 ;
        RECT 6.33 1.625 6.43 1.725 ;
        RECT 6.33 1.395 6.43 1.495 ;
        RECT 6.33 1.165 6.43 1.265 ;
        RECT 6.33 0.935 6.43 1.035 ;
        RECT 6.46 0.65 6.56 0.75 ;
        RECT 6.69 0.65 6.79 0.75 ;
        RECT 6.92 0.65 7.02 0.75 ;
        RECT 7.07 5.035 7.17 5.135 ;
        RECT 7.07 4.805 7.17 4.905 ;
        RECT 7.07 4.575 7.17 4.675 ;
        RECT 7.07 4.345 7.17 4.445 ;
        RECT 7.07 4.115 7.17 4.215 ;
        RECT 7.07 3.885 7.17 3.985 ;
        RECT 7.07 3.445 7.17 3.545 ;
        RECT 7.07 3.215 7.17 3.315 ;
        RECT 7.07 2.985 7.17 3.085 ;
        RECT 7.07 2.755 7.17 2.855 ;
    END
  END VDDSRC
  OBS
    LAYER MET1 ;
      RECT 0.76 1.005 0.9 10.905 ;
      RECT 1.5 1.005 1.64 10.905 ;
      RECT 2.24 1.005 2.38 10.905 ;
      RECT 2.98 1.005 3.12 10.905 ;
      RECT 3.72 1.005 3.86 10.905 ;
      RECT 4.46 1.005 4.6 10.905 ;
      RECT 5.2 1.005 5.34 10.905 ;
      RECT 5.94 1.005 6.08 10.905 ;
      RECT 6.68 1.005 6.82 10.905 ;
      RECT 7.42 1.005 7.56 10.905 ;
      RECT 0.39 0.63 7.56 0.77 ;
      RECT 0.39 0.63 0.53 10.905 ;
      RECT 1.13 0.63 1.27 10.905 ;
      RECT 1.87 0.63 2.01 10.905 ;
      RECT 2.61 0.63 2.75 10.905 ;
      RECT 3.35 0.63 3.49 10.905 ;
      RECT 4.09 0.63 4.23 10.905 ;
      RECT 4.83 0.63 4.97 10.905 ;
      RECT 5.57 0.63 5.71 10.905 ;
      RECT 6.31 0.63 6.45 10.905 ;
      RECT 7.05 0.63 7.19 10.905 ;
  END
END DSIPGX2LPSRCL1
MACRO DSIPGX2LPSRCS1
  CLASS RING ;
  ORIGIN 0 0 ;
  FOREIGN DSIPGX2LPSRCS1 0 0 ;
  SIZE 0.96 BY 11.57 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 0.23 0.96 0.37 ;
      LAYER CUT01 ;
        RECT 0.49 0.255 0.58 0.345 ;
        RECT 0.71 0.255 0.8 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE ANALOG ;
      ANTENNAGATEAREA 1.6 LAYER MET1 ;
      ANTENNAGATEAREA 1.6 LAYER MET2 ;
    ANTENNAMAXCUTCAR 13.125 LAYER CUT01 ;
    SUPPLYSENSITIVITY VDDSRC ;
    GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 0.15 5.38 0.29 11.16 ;
        RECT 0.15 11.02 0.84 11.16 ;
      LAYER MET2 ;
        RECT 0.15 5.38 0.29 6.48 ;
      LAYER CUT12 ;
        RECT 0.17 6.34 0.27 6.44 ;
        RECT 0.17 6.11 0.27 6.21 ;
        RECT 0.17 5.88 0.27 5.98 ;
        RECT 0.17 5.65 0.27 5.75 ;
        RECT 0.17 5.42 0.27 5.52 ;
      LAYER CUT01 ;
        RECT 0.49 11.045 0.58 11.135 ;
        RECT 0.71 11.045 0.8 11.135 ;
    END
  END A
  PIN VDDPD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 0 9.81 0.96 11.25 ;
        RECT 0 8.22 0.96 9.66 ;
        RECT 0 6.63 0.96 8.07 ;
      LAYER CUT12 ;
        RECT 0.78 10.765 0.88 10.865 ;
        RECT 0.78 10.535 0.88 10.635 ;
        RECT 0.78 10.305 0.88 10.405 ;
        RECT 0.78 10.075 0.88 10.175 ;
        RECT 0.78 9.845 0.88 9.945 ;
        RECT 0.78 9.465 0.88 9.565 ;
        RECT 0.78 9.235 0.88 9.335 ;
        RECT 0.78 9.005 0.88 9.105 ;
        RECT 0.78 8.775 0.88 8.875 ;
        RECT 0.78 8.545 0.88 8.645 ;
        RECT 0.78 8.315 0.88 8.415 ;
        RECT 0.78 7.875 0.88 7.975 ;
        RECT 0.78 7.645 0.88 7.745 ;
        RECT 0.78 7.415 0.88 7.515 ;
        RECT 0.78 7.185 0.88 7.285 ;
        RECT 0.78 6.955 0.88 7.055 ;
        RECT 0.78 6.725 0.88 6.825 ;
    END
  END VDDPD
  PIN VDDSRC
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 0 3.79 0.96 5.23 ;
        RECT 0 2.2 0.96 3.64 ;
        RECT 0 0.61 0.96 2.05 ;
      LAYER CUT12 ;
        RECT 0.41 5.035 0.51 5.135 ;
        RECT 0.41 4.805 0.51 4.905 ;
        RECT 0.41 4.575 0.51 4.675 ;
        RECT 0.41 4.345 0.51 4.445 ;
        RECT 0.41 4.115 0.51 4.215 ;
        RECT 0.41 3.885 0.51 3.985 ;
        RECT 0.41 3.445 0.51 3.545 ;
        RECT 0.41 3.215 0.51 3.315 ;
        RECT 0.41 2.985 0.51 3.085 ;
        RECT 0.41 2.755 0.51 2.855 ;
        RECT 0.41 2.525 0.51 2.625 ;
        RECT 0.41 2.295 0.51 2.395 ;
        RECT 0.41 1.855 0.51 1.955 ;
        RECT 0.41 1.625 0.51 1.725 ;
        RECT 0.41 1.395 0.51 1.495 ;
        RECT 0.41 1.165 0.51 1.265 ;
        RECT 0.41 0.935 0.51 1.035 ;
        RECT 0.45 0.65 0.55 0.75 ;
        RECT 0.68 0.65 0.78 0.75 ;
    END
  END VDDSRC
  OBS
    LAYER MET1 ;
      RECT 0.39 0.63 0.84 0.77 ;
      RECT 0.39 0.63 0.53 10.905 ;
      RECT 0.76 1.005 0.9 10.905 ;
  END
END DSIPGX2LPSRCS1
MACRO DSIPGX2LPSRCS2
  CLASS RING ;
  ORIGIN 0 0 ;
  FOREIGN DSIPGX2LPSRCS2 0 0 ;
  SIZE 1.92 BY 11.57 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 0.23 1.92 0.37 ;
      LAYER CUT01 ;
        RECT 0.49 0.255 0.58 0.345 ;
        RECT 0.71 0.255 0.8 0.345 ;
    END
  END VSS
  PIN A
    DIRECTION INPUT ;
    USE ANALOG ;
      ANTENNAGATEAREA 1.6 LAYER MET1 ;
      ANTENNAGATEAREA 1.6 LAYER MET2 ;
    ANTENNAMAXCUTCAR 13.125 LAYER CUT01 ;
    SUPPLYSENSITIVITY VDDSRC ;
    GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 0.15 5.38 0.29 11.16 ;
        RECT 0.15 11.02 0.84 11.16 ;
      LAYER MET2 ;
        RECT 0.15 5.38 0.29 6.48 ;
      LAYER CUT12 ;
        RECT 0.17 6.34 0.27 6.44 ;
        RECT 0.17 6.11 0.27 6.21 ;
        RECT 0.17 5.88 0.27 5.98 ;
        RECT 0.17 5.65 0.27 5.75 ;
        RECT 0.17 5.42 0.27 5.52 ;
      LAYER CUT01 ;
        RECT 0.49 11.045 0.58 11.135 ;
        RECT 0.71 11.045 0.8 11.135 ;
    END
  END A
  PIN VDDPD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 0 9.81 1.92 11.25 ;
        RECT 0 8.22 1.92 9.66 ;
        RECT 0 6.63 1.92 8.07 ;
      LAYER CUT12 ;
        RECT 0.78 10.765 0.88 10.865 ;
        RECT 0.78 10.535 0.88 10.635 ;
        RECT 0.78 10.305 0.88 10.405 ;
        RECT 0.78 10.075 0.88 10.175 ;
        RECT 0.78 9.845 0.88 9.945 ;
        RECT 0.78 9.465 0.88 9.565 ;
        RECT 0.78 9.235 0.88 9.335 ;
        RECT 0.78 9.005 0.88 9.105 ;
        RECT 0.78 8.775 0.88 8.875 ;
        RECT 0.78 8.545 0.88 8.645 ;
        RECT 0.78 8.315 0.88 8.415 ;
        RECT 0.78 7.875 0.88 7.975 ;
        RECT 0.78 7.645 0.88 7.745 ;
        RECT 0.78 7.415 0.88 7.515 ;
        RECT 0.78 7.185 0.88 7.285 ;
        RECT 0.78 6.955 0.88 7.055 ;
        RECT 0.78 6.725 0.88 6.825 ;
    END
  END VDDPD
  PIN VDDSRC
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 0 3.79 1.92 5.23 ;
        RECT 0 2.2 1.92 3.64 ;
        RECT 0 0.61 1.92 2.05 ;
      LAYER CUT12 ;
        RECT 0.41 5.035 0.51 5.135 ;
        RECT 0.41 4.805 0.51 4.905 ;
        RECT 0.41 4.575 0.51 4.675 ;
        RECT 0.41 4.345 0.51 4.445 ;
        RECT 0.41 4.115 0.51 4.215 ;
        RECT 0.41 3.885 0.51 3.985 ;
        RECT 0.41 3.445 0.51 3.545 ;
        RECT 0.41 3.215 0.51 3.315 ;
        RECT 0.41 2.985 0.51 3.085 ;
        RECT 0.41 2.755 0.51 2.855 ;
        RECT 0.41 2.525 0.51 2.625 ;
        RECT 0.41 2.295 0.51 2.395 ;
        RECT 0.41 1.855 0.51 1.955 ;
        RECT 0.41 1.625 0.51 1.725 ;
        RECT 0.41 1.395 0.51 1.495 ;
        RECT 0.41 1.165 0.51 1.265 ;
        RECT 0.41 0.935 0.51 1.035 ;
        RECT 0.45 0.65 0.55 0.75 ;
        RECT 0.68 0.65 0.78 0.75 ;
    END
  END VDDSRC
  OBS
    LAYER MET1 ;
      RECT 0.39 0.63 0.84 0.77 ;
      RECT 0.39 0.63 0.53 10.905 ;
      RECT 0.76 1.005 0.9 10.905 ;
  END
END DSIPGX2LPSRCS2
MACRO DSIPGX2LSPRCS1
  CLASS RING ;
  ORIGIN 0 0 ;
  FOREIGN DSIPGX2LSPRCS1 0 0 ;
  SIZE 0.96 BY 11.57 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 0.23 0.96 0.37 ;
      LAYER CUT01 ;
        RECT 0.49 0.255 0.58 0.345 ;
        RECT 0.71 0.255 0.8 0.345 ;
    END
  END VSS
  PIN VDDPD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 0 9.81 0.96 11.25 ;
        RECT 0 8.22 0.96 9.66 ;
        RECT 0 6.63 0.96 8.07 ;
      LAYER CUT12 ;
        RECT 0.78 10.765 0.88 10.865 ;
        RECT 0.78 10.535 0.88 10.635 ;
        RECT 0.78 10.305 0.88 10.405 ;
        RECT 0.78 10.075 0.88 10.175 ;
        RECT 0.78 9.845 0.88 9.945 ;
        RECT 0.78 9.465 0.88 9.565 ;
        RECT 0.78 9.235 0.88 9.335 ;
        RECT 0.78 9.005 0.88 9.105 ;
        RECT 0.78 8.775 0.88 8.875 ;
        RECT 0.78 8.545 0.88 8.645 ;
        RECT 0.78 8.315 0.88 8.415 ;
        RECT 0.78 7.875 0.88 7.975 ;
        RECT 0.78 7.645 0.88 7.745 ;
        RECT 0.78 7.415 0.88 7.515 ;
        RECT 0.78 7.185 0.88 7.285 ;
        RECT 0.78 6.955 0.88 7.055 ;
        RECT 0.78 6.725 0.88 6.825 ;
    END
  END VDDPD
  PIN VDDSRC
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 0 3.79 0.96 5.23 ;
        RECT 0 2.2 0.96 3.64 ;
        RECT 0 0.61 0.96 2.05 ;
      LAYER CUT12 ;
        RECT 0.41 5.035 0.51 5.135 ;
        RECT 0.41 4.805 0.51 4.905 ;
        RECT 0.41 4.575 0.51 4.675 ;
        RECT 0.41 4.345 0.51 4.445 ;
        RECT 0.41 4.115 0.51 4.215 ;
        RECT 0.41 3.885 0.51 3.985 ;
        RECT 0.41 3.445 0.51 3.545 ;
        RECT 0.41 3.215 0.51 3.315 ;
        RECT 0.41 2.985 0.51 3.085 ;
        RECT 0.41 2.755 0.51 2.855 ;
        RECT 0.41 2.525 0.51 2.625 ;
        RECT 0.41 2.295 0.51 2.395 ;
        RECT 0.41 1.855 0.51 1.955 ;
        RECT 0.41 1.625 0.51 1.725 ;
        RECT 0.41 1.395 0.51 1.495 ;
        RECT 0.41 1.165 0.51 1.265 ;
        RECT 0.41 0.935 0.51 1.035 ;
        RECT 0.45 0.65 0.55 0.75 ;
        RECT 0.68 0.65 0.78 0.75 ;
    END
  END VDDSRC
  OBS
    LAYER MET1 ;
      RECT 0.39 0.63 0.84 0.77 ;
      RECT 0.39 0.63 0.53 5.175 ;
      RECT 0.76 6.685 0.9 10.905 ;
  END
END DSIPGX2LSPRCS1
MACRO DSIPGX2LSPRCS2
  CLASS RING ;
  ORIGIN 0 0 ;
  FOREIGN DSIPGX2LSPRCS2 0 0 ;
  SIZE 1.92 BY 11.57 ;
  SYMMETRY X Y R90 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET1 ;
        RECT 0 0.23 1.92 0.37 ;
      LAYER CUT01 ;
        RECT 0.49 0.255 0.58 0.345 ;
        RECT 0.71 0.255 0.8 0.345 ;
    END
  END VSS
  PIN VDDPD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 0 9.81 1.92 11.25 ;
        RECT 0 8.22 1.92 9.66 ;
        RECT 0 6.63 1.92 8.07 ;
      LAYER CUT12 ;
        RECT 0.78 10.765 0.88 10.865 ;
        RECT 0.78 10.535 0.88 10.635 ;
        RECT 0.78 10.305 0.88 10.405 ;
        RECT 0.78 10.075 0.88 10.175 ;
        RECT 0.78 9.845 0.88 9.945 ;
        RECT 0.78 9.465 0.88 9.565 ;
        RECT 0.78 9.235 0.88 9.335 ;
        RECT 0.78 9.005 0.88 9.105 ;
        RECT 0.78 8.775 0.88 8.875 ;
        RECT 0.78 8.545 0.88 8.645 ;
        RECT 0.78 8.315 0.88 8.415 ;
        RECT 0.78 7.875 0.88 7.975 ;
        RECT 0.78 7.645 0.88 7.745 ;
        RECT 0.78 7.415 0.88 7.515 ;
        RECT 0.78 7.185 0.88 7.285 ;
        RECT 0.78 6.955 0.88 7.055 ;
        RECT 0.78 6.725 0.88 6.825 ;
    END
  END VDDPD
  PIN VDDSRC
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET2 ;
        RECT 0 3.79 1.92 5.23 ;
        RECT 0 2.2 1.92 3.64 ;
        RECT 0 0.61 1.92 2.05 ;
      LAYER CUT12 ;
        RECT 0.41 5.035 0.51 5.135 ;
        RECT 0.41 4.805 0.51 4.905 ;
        RECT 0.41 4.575 0.51 4.675 ;
        RECT 0.41 4.345 0.51 4.445 ;
        RECT 0.41 4.115 0.51 4.215 ;
        RECT 0.41 3.885 0.51 3.985 ;
        RECT 0.41 3.445 0.51 3.545 ;
        RECT 0.41 3.215 0.51 3.315 ;
        RECT 0.41 2.985 0.51 3.085 ;
        RECT 0.41 2.755 0.51 2.855 ;
        RECT 0.41 2.525 0.51 2.625 ;
        RECT 0.41 2.295 0.51 2.395 ;
        RECT 0.41 1.855 0.51 1.955 ;
        RECT 0.41 1.625 0.51 1.725 ;
        RECT 0.41 1.395 0.51 1.495 ;
        RECT 0.41 1.165 0.51 1.265 ;
        RECT 0.41 0.935 0.51 1.035 ;
        RECT 0.45 0.65 0.55 0.75 ;
        RECT 0.68 0.65 0.78 0.75 ;
    END
  END VDDSRC
  OBS
    LAYER MET1 ;
      RECT 0.39 0.63 0.84 0.77 ;
      RECT 0.39 0.63 0.53 5.175 ;
      RECT 0.76 6.685 0.9 10.905 ;
  END
END DSIPGX2LSPRCS2

END LIBRARY
#-------------------------------------------------------------
#-- This Library is the Confidential and Proprietary product
#-- of Fujitsu Limited. Any unauthorized use, reproduction
#-- or transfer of this library is strictly prohibited.
#-- Copyright (c) 2007 by Fujitsu Limited. All Rights Reserved.
#----------------------------------------------------------------
# Revision : 01    2007/06/04
# Comment  : CS202 LVCMOS 7S0G1-12S3G2
# Editer   : FMSL
#----------------------------------------------------------------
VERSION 5.6 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

SITE IOSITE170
  CLASS PAD ;
  SYMMETRY Y ;
  SIZE 0.01 BY 170.00 ;
END IOSITE170

SITE IOSITE141
  CLASS PAD ;
  SYMMETRY Y ;
  SIZE 0.01 BY 141.00 ;
END IOSITE141

SITE IOSITE10
  CLASS PAD ;
  SYMMETRY Y ;
  SIZE 0.01 BY 10.00 ;
END IOSITE10


MACRO IOCB03N00XXA1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB03N00XXA1 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN NC
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END NC
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB03N00XXA1


MACRO IOCB2EBTNH2LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNH2LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNH2LA01


MACRO IOCB2EBTNH4LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNH4LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNH4LA01


MACRO IOCB2EBTNH4NA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNH4NA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNH4NA01


MACRO IOCB2EBTNH6HA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNH6HA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNH6HA01


MACRO IOCB2EBTNH6LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNH6LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNH6LA01


MACRO IOCB2EBTNH8HA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNH8HA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNH8HA01


MACRO IOCB2EBTNH8NA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNH8NA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNH8NA01


MACRO IOCB2EBTNL2LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNL2LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNL2LA01


MACRO IOCB2EBTNL4LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNL4LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNL4LA01


MACRO IOCB2EBTNL4NA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNL4NA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNL4NA01


MACRO IOCB2EBTNL6HA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNL6HA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNL6HA01


MACRO IOCB2EBTNL6LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNL6LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNL6LA01


MACRO IOCB2EBTNL8HA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNL8HA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNL8HA01


MACRO IOCB2EBTNL8NA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNL8NA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNL8NA01


MACRO IOCB2EBTNN2LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNN2LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNN2LA01


MACRO IOCB2EBTNN4LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNN4LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNN4LA01


MACRO IOCB2EBTNN4NA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNN4NA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNN4NA01


MACRO IOCB2EBTNN6HA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNN6HA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNN6HA01


MACRO IOCB2EBTNN6LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNN6LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNN6LA01


MACRO IOCB2EBTNN8HA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNN8HA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNN8HA01


MACRO IOCB2EBTNN8NA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTNN8NA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTNN8NA01


MACRO IOCB2EBTSH2LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSH2LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSH2LA01


MACRO IOCB2EBTSH4LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSH4LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSH4LA01


MACRO IOCB2EBTSH4NA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSH4NA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSH4NA01


MACRO IOCB2EBTSH6HA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSH6HA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSH6HA01


MACRO IOCB2EBTSH6LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSH6LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSH6LA01


MACRO IOCB2EBTSH8HA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSH8HA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSH8HA01


MACRO IOCB2EBTSH8NA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSH8NA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSH8NA01


MACRO IOCB2EBTSL2LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSL2LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSL2LA01


MACRO IOCB2EBTSL4LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSL4LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSL4LA01


MACRO IOCB2EBTSL4NA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSL4NA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSL4NA01


MACRO IOCB2EBTSL6HA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSL6HA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSL6HA01


MACRO IOCB2EBTSL6LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSL6LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSL6LA01


MACRO IOCB2EBTSL8HA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSL8HA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSL8HA01


MACRO IOCB2EBTSL8NA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSL8NA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSL8NA01


MACRO IOCB2EBTSN2LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSN2LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSN2LA01


MACRO IOCB2EBTSN4LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSN4LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSN4LA01


MACRO IOCB2EBTSN4NA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSN4NA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSN4NA01


MACRO IOCB2EBTSN6HA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSN6HA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSN6HA01


MACRO IOCB2EBTSN6LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSN6LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSN6LA01


MACRO IOCB2EBTSN8HA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSN8HA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSN8HA01


MACRO IOCB2EBTSN8NA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EBTSN8NA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EB
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EB
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EBTSN8NA01


MACRO IOCB2EITNHMXA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EITNHMXA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN EA
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDE ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EA
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EITNHMXA01


MACRO IOCB2EITNLMXA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EITNLMXA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN EA
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDE ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EA
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EITNLMXA01


MACRO IOCB2EITNNMXA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EITNNMXA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN EA
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDE ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EA
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EITNNMXA01


MACRO IOCB2EITPDMXA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EITPDMXA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN EA
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EA
  PIN PC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END PC
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EITPDMXA01


MACRO IOCB2EITSHMXA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EITSHMXA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN EA
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDE ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EA
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EITSHMXA01


MACRO IOCB2EITSLMXA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EITSLMXA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN EA
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDE ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EA
  PIN PC
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET2 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET3 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET4 ;
        RECT 23.95 0 24.05 0.5 ;
      LAYER MET5 ;
        RECT 23.95 0 24.05 0.5 ;
    END
  END PC
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EITSLMXA01


MACRO IOCB2EITSNMXA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EITSNMXA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN EA
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDE ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EA
  PIN X
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET2 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET3 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET4 ;
        RECT 35.95 0 36.05 0.5 ;
      LAYER MET5 ;
        RECT 35.95 0 36.05 0.5 ;
    END
  END X
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EITSNMXA01


MACRO IOCB2EOT2X2LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EOT2X2LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN EX
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EX
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EOT2X2LA01


MACRO IOCB2EOT2X4LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EOT2X4LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN EX
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EX
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EOT2X4LA01


MACRO IOCB2EOT2X4NA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EOT2X4NA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN EX
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EX
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EOT2X4NA01


MACRO IOCB2EOT2X6HA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EOT2X6HA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN EX
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EX
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EOT2X6HA01


MACRO IOCB2EOT2X6LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EOT2X6LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN EX
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EX
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EOT2X6LA01


MACRO IOCB2EOT2X8HA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EOT2X8HA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN EX
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EX
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EOT2X8HA01


MACRO IOCB2EOT2X8NA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EOT2X8NA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN EX
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EX
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EOT2X8NA01


MACRO IOCB2EOT3X2LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EOT3X2LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EX
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EX
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EOT3X2LA01


MACRO IOCB2EOT3X4LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EOT3X4LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EX
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EX
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EOT3X4LA01


MACRO IOCB2EOT3X4NA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EOT3X4NA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EX
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EX
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EOT3X4NA01


MACRO IOCB2EOT3X6HA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EOT3X6HA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EX
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EX
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EOT3X6HA01


MACRO IOCB2EOT3X6LA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EOT3X6LA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EX
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EX
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EOT3X6LA01


MACRO IOCB2EOT3X8HA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EOT3X8HA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EX
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EX
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EOT3X8HA01


MACRO IOCB2EOT3X8NA01
  CLASS  PAD ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EOT3X8NA01 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET2 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET3 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET4 ;
        RECT 9.95 0 10.05 0.5 ;
      LAYER MET5 ;
        RECT 9.95 0 10.05 0.5 ;
    END
  END A
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
      SUPPLYSENSITIVITY VDD ;
      GROUNDSENSITIVITY VSS ;
    PORT
      LAYER MET1 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET2 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET3 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET4 ;
        RECT 15.95 0 16.05 0.5 ;
      LAYER MET5 ;
        RECT 15.95 0 16.05 0.5 ;
    END
  END C
  PIN EX
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1 ;
    PORT
      LAYER MET1 ;
        RECT 2 167 38 170 ;
      LAYER MET2 ;
        RECT 2 167 38 170 ;
      LAYER MET3 ;
        RECT 2 167 38 170 ;
      LAYER MET4 ;
        RECT 2 167 38 170 ;
      LAYER MET5 ;
        RECT 2 167 38 170 ;
    END
  END EX
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2EOT3X8NA01


MACRO IOCB2EPD5PI11
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EPD5PI11 0 0 ;
  SIZE 50 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET1 ;
        RECT 7 167 43 170 ;
      LAYER MET2 ;
        RECT 7 167 43 170 ;
      LAYER MET3 ;
        RECT 7 167 43 170 ;
      LAYER MET4 ;
        RECT 7 167 43 170 ;
      LAYER MET5 ;
        RECT 7 167 43 170 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 12.5 50 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 50 19.5 ;
    END
  END VDD
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 50 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 50 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 50 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 50 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 50 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 50 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 50 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 50 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 50 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 50 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 50 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 50 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 50 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 50 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 50 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 50 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 50 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 50 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 50 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 50 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 50 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 50 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 50 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 50 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 50 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 50 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 50 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 50 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 50 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 50 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 50 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 50 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 50 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 50 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 50 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 50 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 50 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 50 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 50 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 50 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 50 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 50 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 50 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 50 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 50 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 50 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 50 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 50 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 50 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 50 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 50 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 50 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 50 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 50 110.6 ;
    END
  END VSS
  OBS
    LAYER MET1 ;
      RECT 0 0 50 170 ;
    LAYER CUT12 ;
      RECT 0 0 50 170 ;
    LAYER MET2 ;
      RECT 0 0 50 170 ;
    LAYER CUT23 ;
      RECT 0 0 50 170 ;
    LAYER MET3 ;
      RECT 0 0 50 170 ;
    LAYER CUT34 ;
      RECT 0 0 50 170 ;
    LAYER MET4 ;
      RECT 0 0 50 170 ;
    LAYER CUT45 ;
      RECT 0 0 50 170 ;
    LAYER MET5 ;
      RECT 0 0 50 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 50.000 2.000 ;
  END
END IOCB2EPD5PI11


MACRO IOCB2EPE5PE11
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EPE5PE11 0 0 ;
  SIZE 50 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 50 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 50 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 50 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 50 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 50 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 50 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 50 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 50 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 50 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 50 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 50 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 50 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 50 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 50 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 50 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 50 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 50 163.5 ;
    END
    PORT
      LAYER MET1 ;
        RECT 7 167 43 170 ;
      LAYER MET2 ;
        RECT 7 167 43 170 ;
      LAYER MET3 ;
        RECT 7 167 43 170 ;
      LAYER MET4 ;
        RECT 7 167 43 170 ;
      LAYER MET5 ;
        RECT 7 167 43 170 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 50 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 50 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 50 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 50 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 50 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 50 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 50 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 50 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 50 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 50 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 50 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 50 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 50 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 50 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 50 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 50 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 50 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 50 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 50 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 50 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 50 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 50 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 50 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 50 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 50 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 50 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 50 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 50 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 50 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 50 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 50 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 50 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 50 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 50 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 50 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 50 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 50 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 50 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 50 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 50 170 ;
    LAYER CUT12 ;
      RECT 0 0 50 170 ;
    LAYER MET2 ;
      RECT 0 0 50 170 ;
    LAYER CUT23 ;
      RECT 0 0 50 170 ;
    LAYER MET3 ;
      RECT 0 0 50 170 ;
    LAYER CUT34 ;
      RECT 0 0 50 170 ;
    LAYER MET4 ;
      RECT 0 0 50 170 ;
    LAYER CUT45 ;
      RECT 0 0 50 170 ;
    LAYER MET5 ;
      RECT 0 0 50 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 50.000 2.000 ;
  END
END IOCB2EPE5PE11


MACRO IOCB2EPG5PB11
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EPG5PB11 0 0 ;
  SIZE 50 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 50 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 50 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 50 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 50 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 50 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 50 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 50 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 50 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 50 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 50 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 50 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 50 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 50 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 50 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 50 151.5 ;
    END
    PORT
      LAYER MET1 ;
        RECT 7 167 43 170 ;
      LAYER MET2 ;
        RECT 7 167 43 170 ;
      LAYER MET3 ;
        RECT 7 167 43 170 ;
      LAYER MET4 ;
        RECT 7 167 43 170 ;
      LAYER MET5 ;
        RECT 7 167 43 170 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 50 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 50 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 50 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 50 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 50 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 50 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 50 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 50 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 50 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 50 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 50 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 50 110.6 ;
    END
  END VSS
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 50 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 50 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 50 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 50 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 50 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 50 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 50 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 50 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 50 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 50 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 50 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 50 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 50 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 50 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 50 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 50 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 50 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 50 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 50 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 50 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 50 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 50 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 50 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 50 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 50 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 50 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 50 139.5 ;
    END
  END VDE
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 50 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 50 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 50 170 ;
    LAYER CUT12 ;
      RECT 0 0 50 170 ;
    LAYER MET2 ;
      RECT 0 0 50 170 ;
    LAYER CUT23 ;
      RECT 0 0 50 170 ;
    LAYER MET3 ;
      RECT 0 0 50 170 ;
    LAYER CUT34 ;
      RECT 0 0 50 170 ;
    LAYER MET4 ;
      RECT 0 0 50 170 ;
    LAYER CUT45 ;
      RECT 0 0 50 170 ;
    LAYER MET5 ;
      RECT 0 0 50 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 50.000 2.000 ;
  END
END IOCB2EPG5PB11


#----------------------------------------------------------------
# Comment  : 07S0G1  CORNER DIVIDER SPACER WIRE PAD
#----------------------------------------------------------------


MACRO ZCGCB2E470XXA1
  CLASS ENDCAP TOPRIGHT ;
  ORIGIN 0 0 ;
  FOREIGN ZCGCB2E470XXA1 0 0 ;
  SIZE 170 BY 170 ;
  SYMMETRY X Y R90 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET5 ;
        RECT 156.5 0 159.5 1 ;
      LAYER MET3 ;
        RECT 158.99 0 161.99 1 ;
      LAYER MET5 ;
        RECT 160.5 0 163.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 152.5 0 155.5 1 ;
      LAYER MET3 ;
        RECT 153.43 0 156.43 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 95.6 0 98.6 1 ;
      LAYER MET5 ;
        RECT 96.5 0 99.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 91.6 0 94.6 1 ;
      LAYER MET5 ;
        RECT 92.5 0 95.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 87.6 0 90.6 1 ;
      LAYER MET5 ;
        RECT 88.5 0 91.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 83.6 0 86.6 1 ;
      LAYER MET5 ;
        RECT 84.5 0 87.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 79.6 0 82.6 1 ;
      LAYER MET5 ;
        RECT 80.5 0 83.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 75.6 0 78.6 1 ;
      LAYER MET5 ;
        RECT 76.5 0 79.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 75.6 1 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 1 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 1 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 1 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 1 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 1 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 1 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 1 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 1 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 1 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 1 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 1 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 1 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 1 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 1 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 1 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 1 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 136.5 0 139.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 128.5 0 131.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 108.5 0 111.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 72.5 0 75.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 64.5 0 67.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 56.5 0 59.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 48.5 0 51.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 40.5 0 43.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 32.5 0 35.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 28.5 0 31.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 1 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 1 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 1 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 1 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 1 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 1 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 1 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 1 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 1 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 1 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET3 ;
        RECT 148.4 0 151.4 1 ;
      LAYER MET5 ;
        RECT 148.5 0 151.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 140.5 0 143.5 1 ;
      LAYER MET3 ;
        RECT 142.84 0 145.84 1 ;
      LAYER MET5 ;
        RECT 144.5 0 147.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 123.6 0 126.6 1 ;
      LAYER MET5 ;
        RECT 124.5 0 127.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 119.6 0 122.6 1 ;
      LAYER MET5 ;
        RECT 120.5 0 123.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 115.6 0 118.6 1 ;
      LAYER MET5 ;
        RECT 116.5 0 119.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 111.6 0 114.6 1 ;
      LAYER MET5 ;
        RECT 112.5 0 115.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 103.6 0 106.6 1 ;
      LAYER MET5 ;
        RECT 104.5 0 107.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 103.6 1 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 1 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 1 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 1 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 1 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 1 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 1 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 1 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 1 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 1 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 1 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 1 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 1 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 1 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 1 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 132.5 0 135.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 100.5 0 103.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 68.5 0 71.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 60.5 0 63.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 52.5 0 55.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 44.5 0 47.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 36.5 0 39.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 24.5 0 27.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 20.5 0 23.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 8.5 0 11.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 4.5 0 7.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 1 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 1 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 1 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 1 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 1 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 1 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 1 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 1 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 1 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 1 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 1 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 107.6 0 110.6 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 1 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET5 ;
        RECT 16.5 0 19.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 12.5 0 15.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 12.5 1 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 1 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 170 170 ;
    LAYER CUT12 ;
      RECT 0 0 170 170 ;
    LAYER MET2 ;
      RECT 0 0 170 170 ;
    LAYER CUT23 ;
      RECT 0 0 170 170 ;
    LAYER MET3 ;
      RECT 0 0 170 170 ;
    LAYER CUT34 ;
      RECT 0 0 170 170 ;
    LAYER MET4 ;
      RECT 0 0 170 170 ;
    LAYER CUT45 ;
      RECT 0 0 170 170 ;
    LAYER MET5 ;
      RECT 0 0 170 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 2.000 2.000 ;
  END
END ZCGCB2E470XXA1


MACRO IOCB2EDA2E4701
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EDA2E4701 0 0 ;
  SIZE 4 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 4 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 4 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 4 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 4 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 4 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 4 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 4 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 4 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 4 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 4 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 4 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 4 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 4 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 4 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 4 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 4 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 4 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 4 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 4 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 4 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 4 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 4 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 4 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 4 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 4 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 4 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 4 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 4 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 4 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 4 170 ;
    LAYER CUT12 ;
      RECT 0 0 4 170 ;
    LAYER MET2 ;
      RECT 0 0 4 170 ;
    LAYER CUT23 ;
      RECT 0 0 4 170 ;
    LAYER MET3 ;
      RECT 0 0 4 170 ;
    LAYER CUT34 ;
      RECT 0 0 4 170 ;
    LAYER MET4 ;
      RECT 0 0 4 170 ;
    LAYER CUT45 ;
      RECT 0 0 4 170 ;
    LAYER MET5 ;
      RECT 0 0 4 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 4.000 2.000 ;
  END
END IOCB2EDA2E4701


MACRO IOCB2EDB2E4701
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EDB2E4701 0 0 ;
  SIZE 4 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  OBS
    LAYER MET1 ;
      RECT 0 0 4 170 ;
    LAYER CUT12 ;
      RECT 0 0 4 170 ;
    LAYER MET2 ;
      RECT 0 0 4 170 ;
    LAYER CUT23 ;
      RECT 0 0 4 170 ;
    LAYER MET3 ;
      RECT 0 0 4 170 ;
    LAYER CUT34 ;
      RECT 0 0 4 170 ;
    LAYER MET4 ;
      RECT 0 0 4 170 ;
    LAYER CUT45 ;
      RECT 0 0 4 170 ;
    LAYER MET5 ;
      RECT 0 0 4 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 4.000 2.000 ;
  END
END IOCB2EDB2E4701


MACRO IOCB2EDC2E4701
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EDC2E4701 0 0 ;
  SIZE 4 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 4 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 4 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 4 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 4 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 4 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 4 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 4 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 4 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 4 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 4 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 4 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 4 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 4 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 4 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 4 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 4 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 4 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 4 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 4 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 4 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 4 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 4 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 4 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 4 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 4 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 4 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 4 110.6 ;
    END
  END VSS
  OBS
    LAYER MET1 ;
      RECT 0 0 4 170 ;
    LAYER CUT12 ;
      RECT 0 0 4 170 ;
    LAYER MET2 ;
      RECT 0 0 4 170 ;
    LAYER CUT23 ;
      RECT 0 0 4 170 ;
    LAYER MET3 ;
      RECT 0 0 4 170 ;
    LAYER CUT34 ;
      RECT 0 0 4 170 ;
    LAYER MET4 ;
      RECT 0 0 4 170 ;
    LAYER CUT45 ;
      RECT 0 0 4 170 ;
    LAYER MET5 ;
      RECT 0 0 4 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 4.000 2.000 ;
  END
END IOCB2EDC2E4701


MACRO IOCB2ES1470A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2ES1470A1 0 0 ;
  SIZE 1 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 1 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 1 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 1 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 1 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 1 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 1 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 1 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 1 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 1 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 1 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 1 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 1 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 1 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 1 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 1 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 1 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 1 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 1 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 1 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 1 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 1 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 1 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 1 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 1 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 1 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 1 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 1 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 1 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 1 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 1 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 1 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 1 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 1 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 1 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 1 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 1 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 1 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 1 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 1 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 1 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 1 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 1 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 1 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 1 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 1 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 1 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 1 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 1 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 1 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 1 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 1 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 1 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 1 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 1 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 1 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 1 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 1 170 ;
    LAYER CUT12 ;
      RECT 0 0 1 170 ;
    LAYER MET2 ;
      RECT 0 0 1 170 ;
    LAYER CUT23 ;
      RECT 0 0 1 170 ;
    LAYER MET3 ;
      RECT 0 0 1 170 ;
    LAYER CUT34 ;
      RECT 0 0 1 170 ;
    LAYER MET4 ;
      RECT 0 0 1 170 ;
    LAYER CUT45 ;
      RECT 0 0 1 170 ;
    LAYER MET5 ;
      RECT 0 0 1 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 1.000 2.000 ;
  END
END IOCB2ES1470A1


MACRO IOCB2ES2470A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2ES2470A1 0 0 ;
  SIZE 2 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 2 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 2 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 2 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 2 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 2 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 2 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 2 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 2 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 2 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 2 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 2 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 2 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 2 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 2 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 2 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 2 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 2 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 2 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 2 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 2 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 2 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 2 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 2 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 2 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 2 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 2 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 2 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 2 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 2 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 2 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 2 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 2 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 2 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 2 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 2 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 2 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 2 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 2 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 2 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 2 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 2 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 2 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 2 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 2 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 2 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 2 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 2 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 2 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 2 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 2 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 2 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 2 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 2 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 2 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 2 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 2 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 2 170 ;
    LAYER CUT12 ;
      RECT 0 0 2 170 ;
    LAYER MET2 ;
      RECT 0 0 2 170 ;
    LAYER CUT23 ;
      RECT 0 0 2 170 ;
    LAYER MET3 ;
      RECT 0 0 2 170 ;
    LAYER CUT34 ;
      RECT 0 0 2 170 ;
    LAYER MET4 ;
      RECT 0 0 2 170 ;
    LAYER CUT45 ;
      RECT 0 0 2 170 ;
    LAYER MET5 ;
      RECT 0 0 2 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 2.000 2.000 ;
  END
END IOCB2ES2470A1


MACRO IOCB2ES5470A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2ES5470A1 0 0 ;
  SIZE 5 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 5 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 5 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 5 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 5 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 5 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 5 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 5 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 5 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 5 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 5 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 5 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 5 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 5 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 5 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 5 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 5 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 5 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 5 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 5 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 5 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 5 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 5 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 5 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 5 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 5 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 5 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 5 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 5 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 5 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 5 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 5 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 5 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 5 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 5 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 5 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 5 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 5 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 5 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 5 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 5 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 5 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 5 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 5 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 5 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 5 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 5 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 5 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 5 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 5 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 5 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 5 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 5 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 5 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 5 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 5 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 5 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 5 170 ;
    LAYER CUT12 ;
      RECT 0 0 5 170 ;
    LAYER MET2 ;
      RECT 0 0 5 170 ;
    LAYER CUT23 ;
      RECT 0 0 5 170 ;
    LAYER MET3 ;
      RECT 0 0 5 170 ;
    LAYER CUT34 ;
      RECT 0 0 5 170 ;
    LAYER MET4 ;
      RECT 0 0 5 170 ;
    LAYER CUT45 ;
      RECT 0 0 5 170 ;
    LAYER MET5 ;
      RECT 0 0 5 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 5.000 2.000 ;
  END
END IOCB2ES5470A1


MACRO IOCB2ESA470A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2ESA470A1 0 0 ;
  SIZE 10 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 10 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 10 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 10 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 10 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 10 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 10 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 10 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 10 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 10 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 10 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 10 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 10 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 10 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 10 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 10 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 10 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 10 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 10 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 10 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 10 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 10 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 10 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 10 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 10 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 10 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 10 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 10 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 10 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 10 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 10 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 10 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 10 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 10 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 10 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 10 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 10 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 10 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 10 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 10 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 10 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 10 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 10 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 10 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 10 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 10 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 10 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 10 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 10 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 10 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 10 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 10 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 10 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 10 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 10 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 10 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 10 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 10 170 ;
    LAYER CUT12 ;
      RECT 0 0 10 170 ;
    LAYER MET2 ;
      RECT 0 0 10 170 ;
    LAYER CUT23 ;
      RECT 0 0 10 170 ;
    LAYER MET3 ;
      RECT 0 0 10 170 ;
    LAYER CUT34 ;
      RECT 0 0 10 170 ;
    LAYER MET4 ;
      RECT 0 0 10 170 ;
    LAYER CUT45 ;
      RECT 0 0 10 170 ;
    LAYER MET5 ;
      RECT 0 0 10 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 10.000 2.000 ;
  END
END IOCB2ESA470A1


MACRO IOCB2ESB470A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2ESB470A1 0 0 ;
  SIZE 0.1 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 0.1 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 0.1 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 0.1 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 0.1 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 0.1 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 0.1 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 0.1 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 0.1 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 0.1 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 0.1 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 0.1 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 0.1 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 0.1 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 0.1 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 0.1 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 0.1 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 0.1 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 0.1 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 0.1 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 0.1 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 0.1 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 0.1 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 0.1 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 0.1 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 0.1 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 0.1 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 0.1 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 0.1 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 0.1 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 0.1 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 0.1 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 0.1 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 0.1 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 0.1 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 0.1 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 0.1 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 0.1 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 0.1 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 0.1 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 0.1 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 0.1 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 0.1 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 0.1 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 0.1 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 0.1 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 0.1 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 0.1 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 0.1 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 0.1 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 0.1 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 0.1 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 0.1 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 0.1 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 0.1 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 0.1 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 0.1 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 0.1 170 ;
    LAYER CUT12 ;
      RECT 0 0 0.1 170 ;
    LAYER MET2 ;
      RECT 0 0 0.1 170 ;
    LAYER CUT23 ;
      RECT 0 0 0.1 170 ;
    LAYER MET3 ;
      RECT 0 0 0.1 170 ;
    LAYER CUT34 ;
      RECT 0 0 0.1 170 ;
    LAYER MET4 ;
      RECT 0 0 0.1 170 ;
    LAYER CUT45 ;
      RECT 0 0 0.1 170 ;
    LAYER MET5 ;
      RECT 0 0 0.1 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 0.100 2.000 ;
  END
END IOCB2ESB470A1


MACRO IOCB2ESD470A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2ESD470A1 0 0 ;
  SIZE 20 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 20 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 20 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 20 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 20 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 20 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 20 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 20 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 20 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 20 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 20 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 20 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 20 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 20 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 20 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 20 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 20 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 20 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 20 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 20 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 20 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 20 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 20 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 20 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 20 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 20 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 20 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 20 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 20 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 20 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 20 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 20 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 20 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 20 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 20 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 20 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 20 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 20 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 20 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 20 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 20 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 20 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 20 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 20 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 20 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 20 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 20 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 20 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 20 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 20 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 20 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 20 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 20 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 20 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 20 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 20 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 20 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 20 170 ;
    LAYER CUT12 ;
      RECT 0 0 20 170 ;
    LAYER MET2 ;
      RECT 0 0 20 170 ;
    LAYER CUT23 ;
      RECT 0 0 20 170 ;
    LAYER MET3 ;
      RECT 0 0 20 170 ;
    LAYER CUT34 ;
      RECT 0 0 20 170 ;
    LAYER MET4 ;
      RECT 0 0 20 170 ;
    LAYER CUT45 ;
      RECT 0 0 20 170 ;
    LAYER MET5 ;
      RECT 0 0 20 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 20.000 2.000 ;
  END
END IOCB2ESD470A1


MACRO IOCB2ESE470A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2ESE470A1 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2ESE470A1


MACRO IOCB2EW3A070A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EW3A070A1 0 0 ;
  SIZE 50 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  OBS
    LAYER CUTG1 ;
      RECT 0 0 50 170 ;
    LAYER METG1 ;
      RECT 0 0 50 170 ;
    LAYER CUTTOP ;
      RECT 0 0 50 170 ;
    LAYER METTOP ;
      RECT 0 0 50 170 ;
      LAYER OVLAP ;
       RECT 0.000 84.000 50.000 86.000 ;
  END
END IOCB2EW3A070A1


MACRO IOCB2EW3A570A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EW3A570A1 0 0 ;
  SIZE 50 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  OBS
    LAYER CUTG1 ;
      RECT 0 0 50 170 ;
    LAYER METG1 ;
      RECT 0 0 50 170 ;
    LAYER CUTTOP ;
      RECT 0 0 50 170 ;
    LAYER METTOP ;
      RECT 0 0 50 170 ;
      LAYER OVLAP ;
       RECT 0.000 84.000 50.000 86.000 ;
  END
END IOCB2EW3A570A1


MACRO IOCB2EWDA070A1
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EWDA070A1 0 0 ;
  SIZE 50 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 14.5 0 20.5 5 ;
      LAYER METTOP ;
        RECT 14.5 0 20.5 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 22 0 28 5 ;
      LAYER METTOP ;
        RECT 22 0 28 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 29.5 0 35.5 5 ;
      LAYER METTOP ;
        RECT 29.5 0 35.5 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 37 0 43 5 ;
      LAYER METTOP ;
        RECT 37 0 43 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 7 0 13 5 ;
      LAYER METTOP ;
        RECT 7 0 13 5 ;
    END
  END VDD
  OBS
    LAYER CUTG1 ;
      RECT 0 0 50 170 ;
    LAYER METG1 ;
      RECT 0 0 50 170 ;
    LAYER CUTTOP ;
      RECT 0 0 50 170 ;
    LAYER METTOP ;
      RECT 0 0 50 170 ;
      LAYER OVLAP ;
       RECT 0.000 84.000 50.000 86.000 ;
  END
END IOCB2EWDA070A1


MACRO IOCB2EWDA570A1
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EWDA570A1 0 0 ;
  SIZE 50 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 14.5 0 20.5 5 ;
      LAYER METTOP ;
        RECT 14.5 0 20.5 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 22 0 28 5 ;
      LAYER METTOP ;
        RECT 22 0 28 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 29.5 0 35.5 5 ;
      LAYER METTOP ;
        RECT 29.5 0 35.5 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 37 0 43 5 ;
      LAYER METTOP ;
        RECT 37 0 43 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 7 0 13 5 ;
      LAYER METTOP ;
        RECT 7 0 13 5 ;
    END
  END VDD
  OBS
    LAYER CUTG1 ;
      RECT 0 0 50 170 ;
    LAYER METG1 ;
      RECT 0 0 50 170 ;
    LAYER CUTTOP ;
      RECT 0 0 50 170 ;
    LAYER METTOP ;
      RECT 0 0 50 170 ;
      LAYER OVLAP ;
       RECT 0.000 84.000 50.000 86.000 ;
  END
END IOCB2EWDA570A1


MACRO IOCB2EWGA070A1
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EWGA070A1 0 0 ;
  SIZE 50 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 14.5 0 20.5 5 ;
      LAYER METTOP ;
        RECT 14.5 0 20.5 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 22 0 28 5 ;
      LAYER METTOP ;
        RECT 22 0 28 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 29.5 0 35.5 5 ;
      LAYER METTOP ;
        RECT 29.5 0 35.5 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 37 0 43 5 ;
      LAYER METTOP ;
        RECT 37 0 43 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 7 0 13 5 ;
      LAYER METTOP ;
        RECT 7 0 13 5 ;
    END
  END VSS
  OBS
    LAYER CUTG1 ;
      RECT 0 0 50 170 ;
    LAYER METG1 ;
      RECT 0 0 50 170 ;
    LAYER CUTTOP ;
      RECT 0 0 50 170 ;
    LAYER METTOP ;
      RECT 0 0 50 170 ;
      LAYER OVLAP ;
       RECT 0.000 84.000 50.000 86.000 ;
  END
END IOCB2EWGA070A1


MACRO IOCB2EWGA570A1
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EWGA570A1 0 0 ;
  SIZE 50 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 14.5 0 20.5 5 ;
      LAYER METTOP ;
        RECT 14.5 0 20.5 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 22 0 28 5 ;
      LAYER METTOP ;
        RECT 22 0 28 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 29.5 0 35.5 5 ;
      LAYER METTOP ;
        RECT 29.5 0 35.5 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 37 0 43 5 ;
      LAYER METTOP ;
        RECT 37 0 43 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG1 ;
        RECT 7 0 13 5 ;
      LAYER METTOP ;
        RECT 7 0 13 5 ;
    END
  END VSS
  OBS
    LAYER CUTG1 ;
      RECT 0 0 50 170 ;
    LAYER METG1 ;
      RECT 0 0 50 170 ;
    LAYER CUTTOP ;
      RECT 0 0 50 170 ;
    LAYER METTOP ;
      RECT 0 0 50 170 ;
      LAYER OVLAP ;
       RECT 0.000 84.000 50.000 86.000 ;
  END
END IOCB2EWGA570A1


MACRO IOCB2EWSA570A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EWSA570A1 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  OBS
    LAYER CUTG1 ;
      RECT 0 0 40 170 ;
    LAYER METG1 ;
      RECT 0 0 40 170 ;
    LAYER CUTTOP ;
      RECT 0 0 40 170 ;
    LAYER METTOP ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 84.000 40.000 86.000 ;
  END
END IOCB2EWSA570A1


MACRO EXTGFCB2E25X70A0
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN EXTGFCB2E25X70A0 0 0 ;
  SIZE 48 BY 141 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE141 ;
  OBS
    LAYER METG1 ;
      RECT 0 0 48 141 ;
    LAYER CUTTOP ;
      RECT 0 0 48 141 ;
    LAYER METTOP ;
      RECT 0 0 48 141 ;
      LAYER OVLAP ;
       RECT 0.000 139.000 48.000 141.000 ;
  END
END EXTGFCB2E25X70A0


#----------------------------------------------------------------
# Comment  : 12S3G2  CORNER DIVIDER SPACER WIRE PAD
#----------------------------------------------------------------

MACRO ZCGCB2E4C0XXA1
  CLASS ENDCAP TOPRIGHT ;
  ORIGIN 0 0 ;
  FOREIGN ZCGCB2E4C0XXA1 0 0 ;
  SIZE 170 BY 170 ;
  SYMMETRY X Y R90 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET5 ;
        RECT 136.5 0 139.5 1 ;
      LAYER MET6 ;
        RECT 136.5 0 139.5 1 ;
      LAYER METG1 ;
        RECT 136.5 0 139.5 1 ;
      LAYER METS1 ;
        RECT 136.5 0 139.5 1 ;
      LAYER METS2 ;
        RECT 136.5 0 139.5 1 ;
      LAYER METS3 ;
        RECT 136.5 0 139.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 128.5 0 131.5 1 ;
      LAYER MET6 ;
        RECT 128.5 0 131.5 1 ;
      LAYER METG1 ;
        RECT 128.5 0 131.5 1 ;
      LAYER METS1 ;
        RECT 128.5 0 131.5 1 ;
      LAYER METS2 ;
        RECT 128.5 0 131.5 1 ;
      LAYER METS3 ;
        RECT 128.5 0 131.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 108.5 0 111.5 1 ;
      LAYER MET6 ;
        RECT 108.5 0 111.5 1 ;
      LAYER METG1 ;
        RECT 108.5 0 111.5 1 ;
      LAYER METS1 ;
        RECT 108.5 0 111.5 1 ;
      LAYER METS2 ;
        RECT 108.5 0 111.5 1 ;
      LAYER METS3 ;
        RECT 108.5 0 111.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 72.5 0 75.5 1 ;
      LAYER MET6 ;
        RECT 72.5 0 75.5 1 ;
      LAYER METG1 ;
        RECT 72.5 0 75.5 1 ;
      LAYER METS1 ;
        RECT 72.5 0 75.5 1 ;
      LAYER METS2 ;
        RECT 72.5 0 75.5 1 ;
      LAYER METS3 ;
        RECT 72.5 0 75.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 64.5 0 67.5 1 ;
      LAYER MET6 ;
        RECT 64.5 0 67.5 1 ;
      LAYER METG1 ;
        RECT 64.5 0 67.5 1 ;
      LAYER METS1 ;
        RECT 64.5 0 67.5 1 ;
      LAYER METS2 ;
        RECT 64.5 0 67.5 1 ;
      LAYER METS3 ;
        RECT 64.5 0 67.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 56.5 0 59.5 1 ;
      LAYER MET6 ;
        RECT 56.5 0 59.5 1 ;
      LAYER METG1 ;
        RECT 56.5 0 59.5 1 ;
      LAYER METS1 ;
        RECT 56.5 0 59.5 1 ;
      LAYER METS2 ;
        RECT 56.5 0 59.5 1 ;
      LAYER METS3 ;
        RECT 56.5 0 59.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 48.5 0 51.5 1 ;
      LAYER MET6 ;
        RECT 48.5 0 51.5 1 ;
      LAYER METG1 ;
        RECT 48.5 0 51.5 1 ;
      LAYER METS1 ;
        RECT 48.5 0 51.5 1 ;
      LAYER METS2 ;
        RECT 48.5 0 51.5 1 ;
      LAYER METS3 ;
        RECT 48.5 0 51.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 40.5 0 43.5 1 ;
      LAYER MET6 ;
        RECT 40.5 0 43.5 1 ;
      LAYER METG1 ;
        RECT 40.5 0 43.5 1 ;
      LAYER METS1 ;
        RECT 40.5 0 43.5 1 ;
      LAYER METS2 ;
        RECT 40.5 0 43.5 1 ;
      LAYER METS3 ;
        RECT 40.5 0 43.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 32.5 0 35.5 1 ;
      LAYER MET6 ;
        RECT 32.5 0 35.5 1 ;
      LAYER METG1 ;
        RECT 32.5 0 35.5 1 ;
      LAYER METS1 ;
        RECT 32.5 0 35.5 1 ;
      LAYER METS2 ;
        RECT 32.5 0 35.5 1 ;
      LAYER METS3 ;
        RECT 32.5 0 35.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 28.5 0 31.5 1 ;
      LAYER MET6 ;
        RECT 28.5 0 31.5 1 ;
      LAYER METG1 ;
        RECT 28.5 0 31.5 1 ;
      LAYER METS1 ;
        RECT 28.5 0 31.5 1 ;
      LAYER METS2 ;
        RECT 28.5 0 31.5 1 ;
      LAYER METS3 ;
        RECT 28.5 0 31.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 28.5 1 31.5 ;
      LAYER MET6 ;
        RECT 0 28.5 1 31.5 ;
      LAYER METG1 ;
        RECT 0 28.5 1 31.5 ;
      LAYER METS1 ;
        RECT 0 28.5 1 31.5 ;
      LAYER METS2 ;
        RECT 0 28.5 1 31.5 ;
      LAYER METS3 ;
        RECT 0 28.5 1 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 1 35.5 ;
      LAYER MET6 ;
        RECT 0 32.5 1 35.5 ;
      LAYER METG1 ;
        RECT 0 32.5 1 35.5 ;
      LAYER METS1 ;
        RECT 0 32.5 1 35.5 ;
      LAYER METS2 ;
        RECT 0 32.5 1 35.5 ;
      LAYER METS3 ;
        RECT 0 32.5 1 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 1 43.5 ;
      LAYER MET6 ;
        RECT 0 40.5 1 43.5 ;
      LAYER METG1 ;
        RECT 0 40.5 1 43.5 ;
      LAYER METS1 ;
        RECT 0 40.5 1 43.5 ;
      LAYER METS2 ;
        RECT 0 40.5 1 43.5 ;
      LAYER METS3 ;
        RECT 0 40.5 1 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 1 51.5 ;
      LAYER MET6 ;
        RECT 0 48.5 1 51.5 ;
      LAYER METG1 ;
        RECT 0 48.5 1 51.5 ;
      LAYER METS1 ;
        RECT 0 48.5 1 51.5 ;
      LAYER METS2 ;
        RECT 0 48.5 1 51.5 ;
      LAYER METS3 ;
        RECT 0 48.5 1 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 1 59.5 ;
      LAYER MET6 ;
        RECT 0 56.5 1 59.5 ;
      LAYER METG1 ;
        RECT 0 56.5 1 59.5 ;
      LAYER METS1 ;
        RECT 0 56.5 1 59.5 ;
      LAYER METS2 ;
        RECT 0 56.5 1 59.5 ;
      LAYER METS3 ;
        RECT 0 56.5 1 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 1 67.5 ;
      LAYER MET6 ;
        RECT 0 64.5 1 67.5 ;
      LAYER METG1 ;
        RECT 0 64.5 1 67.5 ;
      LAYER METS1 ;
        RECT 0 64.5 1 67.5 ;
      LAYER METS2 ;
        RECT 0 64.5 1 67.5 ;
      LAYER METS3 ;
        RECT 0 64.5 1 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 1 75.5 ;
      LAYER MET6 ;
        RECT 0 72.5 1 75.5 ;
      LAYER METG1 ;
        RECT 0 72.5 1 75.5 ;
      LAYER METS1 ;
        RECT 0 72.5 1 75.5 ;
      LAYER METS2 ;
        RECT 0 72.5 1 75.5 ;
      LAYER METS3 ;
        RECT 0 72.5 1 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 1 111.5 ;
      LAYER MET6 ;
        RECT 0 108.5 1 111.5 ;
      LAYER METG1 ;
        RECT 0 108.5 1 111.5 ;
      LAYER METS1 ;
        RECT 0 108.5 1 111.5 ;
      LAYER METS2 ;
        RECT 0 108.5 1 111.5 ;
      LAYER METS3 ;
        RECT 0 108.5 1 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 1 131.5 ;
      LAYER MET6 ;
        RECT 0 128.5 1 131.5 ;
      LAYER METG1 ;
        RECT 0 128.5 1 131.5 ;
      LAYER METS1 ;
        RECT 0 128.5 1 131.5 ;
      LAYER METS2 ;
        RECT 0 128.5 1 131.5 ;
      LAYER METS3 ;
        RECT 0 128.5 1 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 1 139.5 ;
      LAYER MET6 ;
        RECT 0 136.5 1 139.5 ;
      LAYER METG1 ;
        RECT 0 136.5 1 139.5 ;
      LAYER METS1 ;
        RECT 0 136.5 1 139.5 ;
      LAYER METS2 ;
        RECT 0 136.5 1 139.5 ;
      LAYER METS3 ;
        RECT 0 136.5 1 139.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 156.5 0 159.5 1 ;
      LAYER MET6 ;
        RECT 156.5 0 159.5 1 ;
      LAYER METG1 ;
        RECT 156.5 0 159.5 1 ;
      LAYER METS1 ;
        RECT 156.5 0 159.5 1 ;
      LAYER METS2 ;
        RECT 156.5 0 159.5 1 ;
      LAYER METS3 ;
        RECT 156.5 0 159.5 1 ;
      LAYER MET3 ;
        RECT 158.99 0 161.99 1 ;
      LAYER MET5 ;
        RECT 160.5 0 163.5 1 ;
      LAYER MET6 ;
        RECT 160.5 0 163.5 1 ;
      LAYER METG1 ;
        RECT 160.5 0 163.5 1 ;
      LAYER METS1 ;
        RECT 160.5 0 163.5 1 ;
      LAYER METS2 ;
        RECT 160.5 0 163.5 1 ;
      LAYER METS3 ;
        RECT 160.5 0 163.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 152.5 0 155.5 1 ;
      LAYER MET6 ;
        RECT 152.5 0 155.5 1 ;
      LAYER METG1 ;
        RECT 152.5 0 155.5 1 ;
      LAYER METS1 ;
        RECT 152.5 0 155.5 1 ;
      LAYER METS2 ;
        RECT 152.5 0 155.5 1 ;
      LAYER METS3 ;
        RECT 152.5 0 155.5 1 ;
      LAYER MET3 ;
        RECT 153.43 0 156.43 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 95.6 0 98.6 1 ;
      LAYER MET5 ;
        RECT 96.5 0 99.5 1 ;
      LAYER MET6 ;
        RECT 96.5 0 99.5 1 ;
      LAYER METG1 ;
        RECT 96.5 0 99.5 1 ;
      LAYER METS1 ;
        RECT 96.5 0 99.5 1 ;
      LAYER METS2 ;
        RECT 96.5 0 99.5 1 ;
      LAYER METS3 ;
        RECT 96.5 0 99.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 91.6 0 94.6 1 ;
      LAYER MET5 ;
        RECT 92.5 0 95.5 1 ;
      LAYER MET6 ;
        RECT 92.5 0 95.5 1 ;
      LAYER METG1 ;
        RECT 92.5 0 95.5 1 ;
      LAYER METS1 ;
        RECT 92.5 0 95.5 1 ;
      LAYER METS2 ;
        RECT 92.5 0 95.5 1 ;
      LAYER METS3 ;
        RECT 92.5 0 95.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 87.6 0 90.6 1 ;
      LAYER MET5 ;
        RECT 88.5 0 91.5 1 ;
      LAYER MET6 ;
        RECT 88.5 0 91.5 1 ;
      LAYER METG1 ;
        RECT 88.5 0 91.5 1 ;
      LAYER METS1 ;
        RECT 88.5 0 91.5 1 ;
      LAYER METS2 ;
        RECT 88.5 0 91.5 1 ;
      LAYER METS3 ;
        RECT 88.5 0 91.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 83.6 0 86.6 1 ;
      LAYER MET5 ;
        RECT 84.5 0 87.5 1 ;
      LAYER MET6 ;
        RECT 84.5 0 87.5 1 ;
      LAYER METG1 ;
        RECT 84.5 0 87.5 1 ;
      LAYER METS1 ;
        RECT 84.5 0 87.5 1 ;
      LAYER METS2 ;
        RECT 84.5 0 87.5 1 ;
      LAYER METS3 ;
        RECT 84.5 0 87.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 79.6 0 82.6 1 ;
      LAYER MET5 ;
        RECT 80.5 0 83.5 1 ;
      LAYER MET6 ;
        RECT 80.5 0 83.5 1 ;
      LAYER METG1 ;
        RECT 80.5 0 83.5 1 ;
      LAYER METS1 ;
        RECT 80.5 0 83.5 1 ;
      LAYER METS2 ;
        RECT 80.5 0 83.5 1 ;
      LAYER METS3 ;
        RECT 80.5 0 83.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 75.6 0 78.6 1 ;
      LAYER MET5 ;
        RECT 76.5 0 79.5 1 ;
      LAYER MET6 ;
        RECT 76.5 0 79.5 1 ;
      LAYER METG1 ;
        RECT 76.5 0 79.5 1 ;
      LAYER METS1 ;
        RECT 76.5 0 79.5 1 ;
      LAYER METS2 ;
        RECT 76.5 0 79.5 1 ;
      LAYER METS3 ;
        RECT 76.5 0 79.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 75.6 1 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 1 79.5 ;
      LAYER MET6 ;
        RECT 0 76.5 1 79.5 ;
      LAYER METG1 ;
        RECT 0 76.5 1 79.5 ;
      LAYER METS1 ;
        RECT 0 76.5 1 79.5 ;
      LAYER METS2 ;
        RECT 0 76.5 1 79.5 ;
      LAYER METS3 ;
        RECT 0 76.5 1 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 1 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 1 83.5 ;
      LAYER MET6 ;
        RECT 0 80.5 1 83.5 ;
      LAYER METG1 ;
        RECT 0 80.5 1 83.5 ;
      LAYER METS1 ;
        RECT 0 80.5 1 83.5 ;
      LAYER METS2 ;
        RECT 0 80.5 1 83.5 ;
      LAYER METS3 ;
        RECT 0 80.5 1 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 1 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 1 87.5 ;
      LAYER MET6 ;
        RECT 0 84.5 1 87.5 ;
      LAYER METG1 ;
        RECT 0 84.5 1 87.5 ;
      LAYER METS1 ;
        RECT 0 84.5 1 87.5 ;
      LAYER METS2 ;
        RECT 0 84.5 1 87.5 ;
      LAYER METS3 ;
        RECT 0 84.5 1 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 1 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 1 91.5 ;
      LAYER MET6 ;
        RECT 0 88.5 1 91.5 ;
      LAYER METG1 ;
        RECT 0 88.5 1 91.5 ;
      LAYER METS1 ;
        RECT 0 88.5 1 91.5 ;
      LAYER METS2 ;
        RECT 0 88.5 1 91.5 ;
      LAYER METS3 ;
        RECT 0 88.5 1 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 1 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 1 95.5 ;
      LAYER MET6 ;
        RECT 0 92.5 1 95.5 ;
      LAYER METG1 ;
        RECT 0 92.5 1 95.5 ;
      LAYER METS1 ;
        RECT 0 92.5 1 95.5 ;
      LAYER METS2 ;
        RECT 0 92.5 1 95.5 ;
      LAYER METS3 ;
        RECT 0 92.5 1 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 1 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 1 99.5 ;
      LAYER MET6 ;
        RECT 0 96.5 1 99.5 ;
      LAYER METG1 ;
        RECT 0 96.5 1 99.5 ;
      LAYER METS1 ;
        RECT 0 96.5 1 99.5 ;
      LAYER METS2 ;
        RECT 0 96.5 1 99.5 ;
      LAYER METS3 ;
        RECT 0 96.5 1 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 1 155.5 ;
      LAYER MET6 ;
        RECT 0 152.5 1 155.5 ;
      LAYER METG1 ;
        RECT 0 152.5 1 155.5 ;
      LAYER METS1 ;
        RECT 0 152.5 1 155.5 ;
      LAYER METS2 ;
        RECT 0 152.5 1 155.5 ;
      LAYER METS3 ;
        RECT 0 152.5 1 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 1 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 1 159.5 ;
      LAYER MET6 ;
        RECT 0 156.5 1 159.5 ;
      LAYER METG1 ;
        RECT 0 156.5 1 159.5 ;
      LAYER METS1 ;
        RECT 0 156.5 1 159.5 ;
      LAYER METS2 ;
        RECT 0 156.5 1 159.5 ;
      LAYER METS3 ;
        RECT 0 156.5 1 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 1 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 1 163.5 ;
      LAYER MET6 ;
        RECT 0 160.5 1 163.5 ;
      LAYER METG1 ;
        RECT 0 160.5 1 163.5 ;
      LAYER METS1 ;
        RECT 0 160.5 1 163.5 ;
      LAYER METS2 ;
        RECT 0 160.5 1 163.5 ;
      LAYER METS3 ;
        RECT 0 160.5 1 163.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET5 ;
        RECT 132.5 0 135.5 1 ;
      LAYER MET6 ;
        RECT 132.5 0 135.5 1 ;
      LAYER METG1 ;
        RECT 132.5 0 135.5 1 ;
      LAYER METS1 ;
        RECT 132.5 0 135.5 1 ;
      LAYER METS2 ;
        RECT 132.5 0 135.5 1 ;
      LAYER METS3 ;
        RECT 132.5 0 135.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 100.5 0 103.5 1 ;
      LAYER MET6 ;
        RECT 100.5 0 103.5 1 ;
      LAYER METG1 ;
        RECT 100.5 0 103.5 1 ;
      LAYER METS1 ;
        RECT 100.5 0 103.5 1 ;
      LAYER METS2 ;
        RECT 100.5 0 103.5 1 ;
      LAYER METS3 ;
        RECT 100.5 0 103.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 68.5 0 71.5 1 ;
      LAYER MET6 ;
        RECT 68.5 0 71.5 1 ;
      LAYER METG1 ;
        RECT 68.5 0 71.5 1 ;
      LAYER METS1 ;
        RECT 68.5 0 71.5 1 ;
      LAYER METS2 ;
        RECT 68.5 0 71.5 1 ;
      LAYER METS3 ;
        RECT 68.5 0 71.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 60.5 0 63.5 1 ;
      LAYER MET6 ;
        RECT 60.5 0 63.5 1 ;
      LAYER METG1 ;
        RECT 60.5 0 63.5 1 ;
      LAYER METS1 ;
        RECT 60.5 0 63.5 1 ;
      LAYER METS2 ;
        RECT 60.5 0 63.5 1 ;
      LAYER METS3 ;
        RECT 60.5 0 63.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 52.5 0 55.5 1 ;
      LAYER MET6 ;
        RECT 52.5 0 55.5 1 ;
      LAYER METG1 ;
        RECT 52.5 0 55.5 1 ;
      LAYER METS1 ;
        RECT 52.5 0 55.5 1 ;
      LAYER METS2 ;
        RECT 52.5 0 55.5 1 ;
      LAYER METS3 ;
        RECT 52.5 0 55.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 44.5 0 47.5 1 ;
      LAYER MET6 ;
        RECT 44.5 0 47.5 1 ;
      LAYER METG1 ;
        RECT 44.5 0 47.5 1 ;
      LAYER METS1 ;
        RECT 44.5 0 47.5 1 ;
      LAYER METS2 ;
        RECT 44.5 0 47.5 1 ;
      LAYER METS3 ;
        RECT 44.5 0 47.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 36.5 0 39.5 1 ;
      LAYER MET6 ;
        RECT 36.5 0 39.5 1 ;
      LAYER METG1 ;
        RECT 36.5 0 39.5 1 ;
      LAYER METS1 ;
        RECT 36.5 0 39.5 1 ;
      LAYER METS2 ;
        RECT 36.5 0 39.5 1 ;
      LAYER METS3 ;
        RECT 36.5 0 39.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 24.5 0 27.5 1 ;
      LAYER MET6 ;
        RECT 24.5 0 27.5 1 ;
      LAYER METG1 ;
        RECT 24.5 0 27.5 1 ;
      LAYER METS1 ;
        RECT 24.5 0 27.5 1 ;
      LAYER METS2 ;
        RECT 24.5 0 27.5 1 ;
      LAYER METS3 ;
        RECT 24.5 0 27.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 20.5 0 23.5 1 ;
      LAYER MET6 ;
        RECT 20.5 0 23.5 1 ;
      LAYER METG1 ;
        RECT 20.5 0 23.5 1 ;
      LAYER METS1 ;
        RECT 20.5 0 23.5 1 ;
      LAYER METS2 ;
        RECT 20.5 0 23.5 1 ;
      LAYER METS3 ;
        RECT 20.5 0 23.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 8.5 0 11.5 1 ;
      LAYER MET6 ;
        RECT 8.5 0 11.5 1 ;
      LAYER METG1 ;
        RECT 8.5 0 11.5 1 ;
      LAYER METS1 ;
        RECT 8.5 0 11.5 1 ;
      LAYER METS2 ;
        RECT 8.5 0 11.5 1 ;
      LAYER METS3 ;
        RECT 8.5 0 11.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 4.5 0 7.5 1 ;
      LAYER MET6 ;
        RECT 4.5 0 7.5 1 ;
      LAYER METG1 ;
        RECT 4.5 0 7.5 1 ;
      LAYER METS1 ;
        RECT 4.5 0 7.5 1 ;
      LAYER METS2 ;
        RECT 4.5 0 7.5 1 ;
      LAYER METS3 ;
        RECT 4.5 0 7.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 4.5 1 7.5 ;
      LAYER MET6 ;
        RECT 0 4.5 1 7.5 ;
      LAYER METG1 ;
        RECT 0 4.5 1 7.5 ;
      LAYER METS1 ;
        RECT 0 4.5 1 7.5 ;
      LAYER METS2 ;
        RECT 0 4.5 1 7.5 ;
      LAYER METS3 ;
        RECT 0 4.5 1 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 1 11.5 ;
      LAYER MET6 ;
        RECT 0 8.5 1 11.5 ;
      LAYER METG1 ;
        RECT 0 8.5 1 11.5 ;
      LAYER METS1 ;
        RECT 0 8.5 1 11.5 ;
      LAYER METS2 ;
        RECT 0 8.5 1 11.5 ;
      LAYER METS3 ;
        RECT 0 8.5 1 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 1 23.5 ;
      LAYER MET6 ;
        RECT 0 20.5 1 23.5 ;
      LAYER METG1 ;
        RECT 0 20.5 1 23.5 ;
      LAYER METS1 ;
        RECT 0 20.5 1 23.5 ;
      LAYER METS2 ;
        RECT 0 20.5 1 23.5 ;
      LAYER METS3 ;
        RECT 0 20.5 1 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 1 27.5 ;
      LAYER MET6 ;
        RECT 0 24.5 1 27.5 ;
      LAYER METG1 ;
        RECT 0 24.5 1 27.5 ;
      LAYER METS1 ;
        RECT 0 24.5 1 27.5 ;
      LAYER METS2 ;
        RECT 0 24.5 1 27.5 ;
      LAYER METS3 ;
        RECT 0 24.5 1 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 1 39.5 ;
      LAYER MET6 ;
        RECT 0 36.5 1 39.5 ;
      LAYER METG1 ;
        RECT 0 36.5 1 39.5 ;
      LAYER METS1 ;
        RECT 0 36.5 1 39.5 ;
      LAYER METS2 ;
        RECT 0 36.5 1 39.5 ;
      LAYER METS3 ;
        RECT 0 36.5 1 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 1 47.5 ;
      LAYER MET6 ;
        RECT 0 44.5 1 47.5 ;
      LAYER METG1 ;
        RECT 0 44.5 1 47.5 ;
      LAYER METS1 ;
        RECT 0 44.5 1 47.5 ;
      LAYER METS2 ;
        RECT 0 44.5 1 47.5 ;
      LAYER METS3 ;
        RECT 0 44.5 1 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 1 55.5 ;
      LAYER MET6 ;
        RECT 0 52.5 1 55.5 ;
      LAYER METG1 ;
        RECT 0 52.5 1 55.5 ;
      LAYER METS1 ;
        RECT 0 52.5 1 55.5 ;
      LAYER METS2 ;
        RECT 0 52.5 1 55.5 ;
      LAYER METS3 ;
        RECT 0 52.5 1 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 1 63.5 ;
      LAYER MET6 ;
        RECT 0 60.5 1 63.5 ;
      LAYER METG1 ;
        RECT 0 60.5 1 63.5 ;
      LAYER METS1 ;
        RECT 0 60.5 1 63.5 ;
      LAYER METS2 ;
        RECT 0 60.5 1 63.5 ;
      LAYER METS3 ;
        RECT 0 60.5 1 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 1 71.5 ;
      LAYER MET6 ;
        RECT 0 68.5 1 71.5 ;
      LAYER METG1 ;
        RECT 0 68.5 1 71.5 ;
      LAYER METS1 ;
        RECT 0 68.5 1 71.5 ;
      LAYER METS2 ;
        RECT 0 68.5 1 71.5 ;
      LAYER METS3 ;
        RECT 0 68.5 1 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 1 103.5 ;
      LAYER MET6 ;
        RECT 0 100.5 1 103.5 ;
      LAYER METG1 ;
        RECT 0 100.5 1 103.5 ;
      LAYER METS1 ;
        RECT 0 100.5 1 103.5 ;
      LAYER METS2 ;
        RECT 0 100.5 1 103.5 ;
      LAYER METS3 ;
        RECT 0 100.5 1 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 1 135.5 ;
      LAYER MET6 ;
        RECT 0 132.5 1 135.5 ;
      LAYER METG1 ;
        RECT 0 132.5 1 135.5 ;
      LAYER METS1 ;
        RECT 0 132.5 1 135.5 ;
      LAYER METS2 ;
        RECT 0 132.5 1 135.5 ;
      LAYER METS3 ;
        RECT 0 132.5 1 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 148.4 0 151.4 1 ;
      LAYER MET5 ;
        RECT 148.5 0 151.5 1 ;
      LAYER MET6 ;
        RECT 148.5 0 151.5 1 ;
      LAYER METG1 ;
        RECT 148.5 0 151.5 1 ;
      LAYER METS1 ;
        RECT 148.5 0 151.5 1 ;
      LAYER METS2 ;
        RECT 148.5 0 151.5 1 ;
      LAYER METS3 ;
        RECT 148.5 0 151.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 140.5 0 143.5 1 ;
      LAYER MET6 ;
        RECT 140.5 0 143.5 1 ;
      LAYER METG1 ;
        RECT 140.5 0 143.5 1 ;
      LAYER METS1 ;
        RECT 140.5 0 143.5 1 ;
      LAYER METS2 ;
        RECT 140.5 0 143.5 1 ;
      LAYER METS3 ;
        RECT 140.5 0 143.5 1 ;
      LAYER MET3 ;
        RECT 142.84 0 145.84 1 ;
      LAYER MET5 ;
        RECT 144.5 0 147.5 1 ;
      LAYER MET6 ;
        RECT 144.5 0 147.5 1 ;
      LAYER METG1 ;
        RECT 144.5 0 147.5 1 ;
      LAYER METS1 ;
        RECT 144.5 0 147.5 1 ;
      LAYER METS2 ;
        RECT 144.5 0 147.5 1 ;
      LAYER METS3 ;
        RECT 144.5 0 147.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 123.6 0 126.6 1 ;
      LAYER MET5 ;
        RECT 124.5 0 127.5 1 ;
      LAYER MET6 ;
        RECT 124.5 0 127.5 1 ;
      LAYER METG1 ;
        RECT 124.5 0 127.5 1 ;
      LAYER METS1 ;
        RECT 124.5 0 127.5 1 ;
      LAYER METS2 ;
        RECT 124.5 0 127.5 1 ;
      LAYER METS3 ;
        RECT 124.5 0 127.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 119.6 0 122.6 1 ;
      LAYER MET5 ;
        RECT 120.5 0 123.5 1 ;
      LAYER MET6 ;
        RECT 120.5 0 123.5 1 ;
      LAYER METG1 ;
        RECT 120.5 0 123.5 1 ;
      LAYER METS1 ;
        RECT 120.5 0 123.5 1 ;
      LAYER METS2 ;
        RECT 120.5 0 123.5 1 ;
      LAYER METS3 ;
        RECT 120.5 0 123.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 115.6 0 118.6 1 ;
      LAYER MET5 ;
        RECT 116.5 0 119.5 1 ;
      LAYER MET6 ;
        RECT 116.5 0 119.5 1 ;
      LAYER METG1 ;
        RECT 116.5 0 119.5 1 ;
      LAYER METS1 ;
        RECT 116.5 0 119.5 1 ;
      LAYER METS2 ;
        RECT 116.5 0 119.5 1 ;
      LAYER METS3 ;
        RECT 116.5 0 119.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 111.6 0 114.6 1 ;
      LAYER MET5 ;
        RECT 112.5 0 115.5 1 ;
      LAYER MET6 ;
        RECT 112.5 0 115.5 1 ;
      LAYER METG1 ;
        RECT 112.5 0 115.5 1 ;
      LAYER METS1 ;
        RECT 112.5 0 115.5 1 ;
      LAYER METS2 ;
        RECT 112.5 0 115.5 1 ;
      LAYER METS3 ;
        RECT 112.5 0 115.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 103.6 0 106.6 1 ;
      LAYER MET5 ;
        RECT 104.5 0 107.5 1 ;
      LAYER MET6 ;
        RECT 104.5 0 107.5 1 ;
      LAYER METG1 ;
        RECT 104.5 0 107.5 1 ;
      LAYER METS1 ;
        RECT 104.5 0 107.5 1 ;
      LAYER METS2 ;
        RECT 104.5 0 107.5 1 ;
      LAYER METS3 ;
        RECT 104.5 0 107.5 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 103.6 1 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 1 107.5 ;
      LAYER MET6 ;
        RECT 0 104.5 1 107.5 ;
      LAYER METG1 ;
        RECT 0 104.5 1 107.5 ;
      LAYER METS1 ;
        RECT 0 104.5 1 107.5 ;
      LAYER METS2 ;
        RECT 0 104.5 1 107.5 ;
      LAYER METS3 ;
        RECT 0 104.5 1 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 1 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 1 115.5 ;
      LAYER MET6 ;
        RECT 0 112.5 1 115.5 ;
      LAYER METG1 ;
        RECT 0 112.5 1 115.5 ;
      LAYER METS1 ;
        RECT 0 112.5 1 115.5 ;
      LAYER METS2 ;
        RECT 0 112.5 1 115.5 ;
      LAYER METS3 ;
        RECT 0 112.5 1 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 1 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 1 119.5 ;
      LAYER MET6 ;
        RECT 0 116.5 1 119.5 ;
      LAYER METG1 ;
        RECT 0 116.5 1 119.5 ;
      LAYER METS1 ;
        RECT 0 116.5 1 119.5 ;
      LAYER METS2 ;
        RECT 0 116.5 1 119.5 ;
      LAYER METS3 ;
        RECT 0 116.5 1 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 1 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 1 123.5 ;
      LAYER MET6 ;
        RECT 0 120.5 1 123.5 ;
      LAYER METG1 ;
        RECT 0 120.5 1 123.5 ;
      LAYER METS1 ;
        RECT 0 120.5 1 123.5 ;
      LAYER METS2 ;
        RECT 0 120.5 1 123.5 ;
      LAYER METS3 ;
        RECT 0 120.5 1 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 1 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 1 127.5 ;
      LAYER MET6 ;
        RECT 0 124.5 1 127.5 ;
      LAYER METG1 ;
        RECT 0 124.5 1 127.5 ;
      LAYER METS1 ;
        RECT 0 124.5 1 127.5 ;
      LAYER METS2 ;
        RECT 0 124.5 1 127.5 ;
      LAYER METS3 ;
        RECT 0 124.5 1 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 1 143.5 ;
      LAYER MET6 ;
        RECT 0 140.5 1 143.5 ;
      LAYER METG1 ;
        RECT 0 140.5 1 143.5 ;
      LAYER METS1 ;
        RECT 0 140.5 1 143.5 ;
      LAYER METS2 ;
        RECT 0 140.5 1 143.5 ;
      LAYER METS3 ;
        RECT 0 140.5 1 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 1 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 1 147.5 ;
      LAYER MET6 ;
        RECT 0 144.5 1 147.5 ;
      LAYER METG1 ;
        RECT 0 144.5 1 147.5 ;
      LAYER METS1 ;
        RECT 0 144.5 1 147.5 ;
      LAYER METS2 ;
        RECT 0 144.5 1 147.5 ;
      LAYER METS3 ;
        RECT 0 144.5 1 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 1 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 1 151.5 ;
      LAYER MET6 ;
        RECT 0 148.5 1 151.5 ;
      LAYER METG1 ;
        RECT 0 148.5 1 151.5 ;
      LAYER METS1 ;
        RECT 0 148.5 1 151.5 ;
      LAYER METS2 ;
        RECT 0 148.5 1 151.5 ;
      LAYER METS3 ;
        RECT 0 148.5 1 151.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 107.6 0 110.6 1 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 1 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER MET5 ;
        RECT 16.5 0 19.5 1 ;
      LAYER MET6 ;
        RECT 16.5 0 19.5 1 ;
      LAYER METG1 ;
        RECT 16.5 0 19.5 1 ;
      LAYER METS1 ;
        RECT 16.5 0 19.5 1 ;
      LAYER METS2 ;
        RECT 16.5 0 19.5 1 ;
      LAYER METS3 ;
        RECT 16.5 0 19.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 12.5 0 15.5 1 ;
      LAYER MET6 ;
        RECT 12.5 0 15.5 1 ;
      LAYER METG1 ;
        RECT 12.5 0 15.5 1 ;
      LAYER METS1 ;
        RECT 12.5 0 15.5 1 ;
      LAYER METS2 ;
        RECT 12.5 0 15.5 1 ;
      LAYER METS3 ;
        RECT 12.5 0 15.5 1 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 12.5 1 15.5 ;
      LAYER MET6 ;
        RECT 0 12.5 1 15.5 ;
      LAYER METG1 ;
        RECT 0 12.5 1 15.5 ;
      LAYER METS1 ;
        RECT 0 12.5 1 15.5 ;
      LAYER METS2 ;
        RECT 0 12.5 1 15.5 ;
      LAYER METS3 ;
        RECT 0 12.5 1 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 1 19.5 ;
      LAYER MET6 ;
        RECT 0 16.5 1 19.5 ;
      LAYER METG1 ;
        RECT 0 16.5 1 19.5 ;
      LAYER METS1 ;
        RECT 0 16.5 1 19.5 ;
      LAYER METS2 ;
        RECT 0 16.5 1 19.5 ;
      LAYER METS3 ;
        RECT 0 16.5 1 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 170 170 ;
    LAYER CUT12 ;
      RECT 0 0 170 170 ;
    LAYER MET2 ;
      RECT 0 0 170 170 ;
    LAYER CUT23 ;
      RECT 0 0 170 170 ;
    LAYER MET3 ;
      RECT 0 0 170 170 ;
    LAYER CUT34 ;
      RECT 0 0 170 170 ;
    LAYER MET4 ;
      RECT 0 0 170 170 ;
    LAYER CUT45 ;
      RECT 0 0 170 170 ;
    LAYER MET5 ;
      RECT 0 0 170 170 ;
    LAYER CUT56 ;
      RECT 0 0 170 170 ;
    LAYER MET6 ;
      RECT 0 0 170 170 ;
    LAYER CUTS1 ;
      RECT 0 0 170 170 ;
    LAYER METS1 ;
      RECT 0 0 170 170 ;
    LAYER CUTS2 ;
      RECT 0 0 170 170 ;
    LAYER METS2 ;
      RECT 0 0 170 170 ;
    LAYER CUTS3 ;
      RECT 0 0 170 170 ;
    LAYER METS3 ;
      RECT 0 0 170 170 ;
    LAYER CUTG1 ;
      RECT 0 0 170 170 ;
    LAYER METG1 ;
      RECT 0 0 170 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 2.000 2.000 ;
  END
END ZCGCB2E4C0XXA1


MACRO IOCB2EDA2E4C01
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EDA2E4C01 0 0 ;
  SIZE 4 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 4.5 4 7.5 ;
      LAYER MET6 ;
        RECT 0 4.5 4 7.5 ;
      LAYER METG1 ;
        RECT 0 4.5 4 7.5 ;
      LAYER METS1 ;
        RECT 0 4.5 4 7.5 ;
      LAYER METS2 ;
        RECT 0 4.5 4 7.5 ;
      LAYER METS3 ;
        RECT 0 4.5 4 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 4 11.5 ;
      LAYER MET6 ;
        RECT 0 8.5 4 11.5 ;
      LAYER METG1 ;
        RECT 0 8.5 4 11.5 ;
      LAYER METS1 ;
        RECT 0 8.5 4 11.5 ;
      LAYER METS2 ;
        RECT 0 8.5 4 11.5 ;
      LAYER METS3 ;
        RECT 0 8.5 4 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 4 23.5 ;
      LAYER MET6 ;
        RECT 0 20.5 4 23.5 ;
      LAYER METG1 ;
        RECT 0 20.5 4 23.5 ;
      LAYER METS1 ;
        RECT 0 20.5 4 23.5 ;
      LAYER METS2 ;
        RECT 0 20.5 4 23.5 ;
      LAYER METS3 ;
        RECT 0 20.5 4 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 4 27.5 ;
      LAYER MET6 ;
        RECT 0 24.5 4 27.5 ;
      LAYER METG1 ;
        RECT 0 24.5 4 27.5 ;
      LAYER METS1 ;
        RECT 0 24.5 4 27.5 ;
      LAYER METS2 ;
        RECT 0 24.5 4 27.5 ;
      LAYER METS3 ;
        RECT 0 24.5 4 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 4 39.5 ;
      LAYER MET6 ;
        RECT 0 36.5 4 39.5 ;
      LAYER METG1 ;
        RECT 0 36.5 4 39.5 ;
      LAYER METS1 ;
        RECT 0 36.5 4 39.5 ;
      LAYER METS2 ;
        RECT 0 36.5 4 39.5 ;
      LAYER METS3 ;
        RECT 0 36.5 4 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 4 47.5 ;
      LAYER MET6 ;
        RECT 0 44.5 4 47.5 ;
      LAYER METG1 ;
        RECT 0 44.5 4 47.5 ;
      LAYER METS1 ;
        RECT 0 44.5 4 47.5 ;
      LAYER METS2 ;
        RECT 0 44.5 4 47.5 ;
      LAYER METS3 ;
        RECT 0 44.5 4 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 4 55.5 ;
      LAYER MET6 ;
        RECT 0 52.5 4 55.5 ;
      LAYER METG1 ;
        RECT 0 52.5 4 55.5 ;
      LAYER METS1 ;
        RECT 0 52.5 4 55.5 ;
      LAYER METS2 ;
        RECT 0 52.5 4 55.5 ;
      LAYER METS3 ;
        RECT 0 52.5 4 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 4 63.5 ;
      LAYER MET6 ;
        RECT 0 60.5 4 63.5 ;
      LAYER METG1 ;
        RECT 0 60.5 4 63.5 ;
      LAYER METS1 ;
        RECT 0 60.5 4 63.5 ;
      LAYER METS2 ;
        RECT 0 60.5 4 63.5 ;
      LAYER METS3 ;
        RECT 0 60.5 4 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 4 71.5 ;
      LAYER MET6 ;
        RECT 0 68.5 4 71.5 ;
      LAYER METG1 ;
        RECT 0 68.5 4 71.5 ;
      LAYER METS1 ;
        RECT 0 68.5 4 71.5 ;
      LAYER METS2 ;
        RECT 0 68.5 4 71.5 ;
      LAYER METS3 ;
        RECT 0 68.5 4 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 4 103.5 ;
      LAYER MET6 ;
        RECT 0 100.5 4 103.5 ;
      LAYER METG1 ;
        RECT 0 100.5 4 103.5 ;
      LAYER METS1 ;
        RECT 0 100.5 4 103.5 ;
      LAYER METS2 ;
        RECT 0 100.5 4 103.5 ;
      LAYER METS3 ;
        RECT 0 100.5 4 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 4 135.5 ;
      LAYER MET6 ;
        RECT 0 132.5 4 135.5 ;
      LAYER METG1 ;
        RECT 0 132.5 4 135.5 ;
      LAYER METS1 ;
        RECT 0 132.5 4 135.5 ;
      LAYER METS2 ;
        RECT 0 132.5 4 135.5 ;
      LAYER METS3 ;
        RECT 0 132.5 4 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 103.6 4 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 4 107.5 ;
      LAYER MET6 ;
        RECT 0 104.5 4 107.5 ;
      LAYER METG1 ;
        RECT 0 104.5 4 107.5 ;
      LAYER METS1 ;
        RECT 0 104.5 4 107.5 ;
      LAYER METS2 ;
        RECT 0 104.5 4 107.5 ;
      LAYER METS3 ;
        RECT 0 104.5 4 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 4 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 4 115.5 ;
      LAYER MET6 ;
        RECT 0 112.5 4 115.5 ;
      LAYER METG1 ;
        RECT 0 112.5 4 115.5 ;
      LAYER METS1 ;
        RECT 0 112.5 4 115.5 ;
      LAYER METS2 ;
        RECT 0 112.5 4 115.5 ;
      LAYER METS3 ;
        RECT 0 112.5 4 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 4 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 4 119.5 ;
      LAYER MET6 ;
        RECT 0 116.5 4 119.5 ;
      LAYER METG1 ;
        RECT 0 116.5 4 119.5 ;
      LAYER METS1 ;
        RECT 0 116.5 4 119.5 ;
      LAYER METS2 ;
        RECT 0 116.5 4 119.5 ;
      LAYER METS3 ;
        RECT 0 116.5 4 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 4 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 4 123.5 ;
      LAYER MET6 ;
        RECT 0 120.5 4 123.5 ;
      LAYER METG1 ;
        RECT 0 120.5 4 123.5 ;
      LAYER METS1 ;
        RECT 0 120.5 4 123.5 ;
      LAYER METS2 ;
        RECT 0 120.5 4 123.5 ;
      LAYER METS3 ;
        RECT 0 120.5 4 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 4 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 4 127.5 ;
      LAYER MET6 ;
        RECT 0 124.5 4 127.5 ;
      LAYER METG1 ;
        RECT 0 124.5 4 127.5 ;
      LAYER METS1 ;
        RECT 0 124.5 4 127.5 ;
      LAYER METS2 ;
        RECT 0 124.5 4 127.5 ;
      LAYER METS3 ;
        RECT 0 124.5 4 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 4 143.5 ;
      LAYER MET6 ;
        RECT 0 140.5 4 143.5 ;
      LAYER METG1 ;
        RECT 0 140.5 4 143.5 ;
      LAYER METS1 ;
        RECT 0 140.5 4 143.5 ;
      LAYER METS2 ;
        RECT 0 140.5 4 143.5 ;
      LAYER METS3 ;
        RECT 0 140.5 4 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 4 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 4 147.5 ;
      LAYER MET6 ;
        RECT 0 144.5 4 147.5 ;
      LAYER METG1 ;
        RECT 0 144.5 4 147.5 ;
      LAYER METS1 ;
        RECT 0 144.5 4 147.5 ;
      LAYER METS2 ;
        RECT 0 144.5 4 147.5 ;
      LAYER METS3 ;
        RECT 0 144.5 4 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 4 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 4 151.5 ;
      LAYER MET6 ;
        RECT 0 148.5 4 151.5 ;
      LAYER METG1 ;
        RECT 0 148.5 4 151.5 ;
      LAYER METS1 ;
        RECT 0 148.5 4 151.5 ;
      LAYER METS2 ;
        RECT 0 148.5 4 151.5 ;
      LAYER METS3 ;
        RECT 0 148.5 4 151.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 4 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 4 15.5 ;
      LAYER MET6 ;
        RECT 0 12.5 4 15.5 ;
      LAYER METG1 ;
        RECT 0 12.5 4 15.5 ;
      LAYER METS1 ;
        RECT 0 12.5 4 15.5 ;
      LAYER METS2 ;
        RECT 0 12.5 4 15.5 ;
      LAYER METS3 ;
        RECT 0 12.5 4 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 4 19.5 ;
      LAYER MET6 ;
        RECT 0 16.5 4 19.5 ;
      LAYER METG1 ;
        RECT 0 16.5 4 19.5 ;
      LAYER METS1 ;
        RECT 0 16.5 4 19.5 ;
      LAYER METS2 ;
        RECT 0 16.5 4 19.5 ;
      LAYER METS3 ;
        RECT 0 16.5 4 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 4 170 ;
    LAYER CUT12 ;
      RECT 0 0 4 170 ;
    LAYER MET2 ;
      RECT 0 0 4 170 ;
    LAYER CUT23 ;
      RECT 0 0 4 170 ;
    LAYER MET3 ;
      RECT 0 0 4 170 ;
    LAYER CUT34 ;
      RECT 0 0 4 170 ;
    LAYER MET4 ;
      RECT 0 0 4 170 ;
    LAYER CUT45 ;
      RECT 0 0 4 170 ;
    LAYER MET5 ;
      RECT 0 0 4 170 ;
    LAYER CUT56 ;
      RECT 0 0 4 170 ;
    LAYER MET6 ;
      RECT 0 0 4 170 ;
    LAYER CUTS1 ;
      RECT 0 0 4 170 ;
    LAYER METS1 ;
      RECT 0 0 4 170 ;
    LAYER CUTS2 ;
      RECT 0 0 4 170 ;
    LAYER METS2 ;
      RECT 0 0 4 170 ;
    LAYER CUTS3 ;
      RECT 0 0 4 170 ;
    LAYER METS3 ;
      RECT 0 0 4 170 ;
    LAYER CUTG1 ;
      RECT 0 0 4 170 ;
    LAYER METG1 ;
      RECT 0 0 4 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 4.000 2.000 ;
  END
END IOCB2EDA2E4C01


MACRO IOCB2EDB2E4C01
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EDB2E4C01 0 0 ;
  SIZE 4 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  OBS
    LAYER MET1 ;
      RECT 0 0 4 170 ;
    LAYER CUT12 ;
      RECT 0 0 4 170 ;
    LAYER MET2 ;
      RECT 0 0 4 170 ;
    LAYER CUT23 ;
      RECT 0 0 4 170 ;
    LAYER MET3 ;
      RECT 0 0 4 170 ;
    LAYER CUT34 ;
      RECT 0 0 4 170 ;
    LAYER MET4 ;
      RECT 0 0 4 170 ;
    LAYER CUT45 ;
      RECT 0 0 4 170 ;
    LAYER MET5 ;
      RECT 0 0 4 170 ;
    LAYER CUT56 ;
      RECT 0 0 4 170 ;
    LAYER MET6 ;
      RECT 0 0 4 170 ;
    LAYER CUTS1 ;
      RECT 0 0 4 170 ;
    LAYER METS1 ;
      RECT 0 0 4 170 ;
    LAYER CUTS2 ;
      RECT 0 0 4 170 ;
    LAYER METS2 ;
      RECT 0 0 4 170 ;
    LAYER CUTS3 ;
      RECT 0 0 4 170 ;
    LAYER METS3 ;
      RECT 0 0 4 170 ;
    LAYER CUTG1 ;
      RECT 0 0 4 170 ;
    LAYER METG1 ;
      RECT 0 0 4 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 4.000 2.000 ;
  END
END IOCB2EDB2E4C01


MACRO IOCB2EDC2E4C01
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EDC2E4C01 0 0 ;
  SIZE 4 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 4.5 4 7.5 ;
      LAYER MET6 ;
        RECT 0 4.5 4 7.5 ;
      LAYER METG1 ;
        RECT 0 4.5 4 7.5 ;
      LAYER METS1 ;
        RECT 0 4.5 4 7.5 ;
      LAYER METS2 ;
        RECT 0 4.5 4 7.5 ;
      LAYER METS3 ;
        RECT 0 4.5 4 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 4 11.5 ;
      LAYER MET6 ;
        RECT 0 8.5 4 11.5 ;
      LAYER METG1 ;
        RECT 0 8.5 4 11.5 ;
      LAYER METS1 ;
        RECT 0 8.5 4 11.5 ;
      LAYER METS2 ;
        RECT 0 8.5 4 11.5 ;
      LAYER METS3 ;
        RECT 0 8.5 4 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 4 23.5 ;
      LAYER MET6 ;
        RECT 0 20.5 4 23.5 ;
      LAYER METG1 ;
        RECT 0 20.5 4 23.5 ;
      LAYER METS1 ;
        RECT 0 20.5 4 23.5 ;
      LAYER METS2 ;
        RECT 0 20.5 4 23.5 ;
      LAYER METS3 ;
        RECT 0 20.5 4 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 4 27.5 ;
      LAYER MET6 ;
        RECT 0 24.5 4 27.5 ;
      LAYER METG1 ;
        RECT 0 24.5 4 27.5 ;
      LAYER METS1 ;
        RECT 0 24.5 4 27.5 ;
      LAYER METS2 ;
        RECT 0 24.5 4 27.5 ;
      LAYER METS3 ;
        RECT 0 24.5 4 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 4 39.5 ;
      LAYER MET6 ;
        RECT 0 36.5 4 39.5 ;
      LAYER METG1 ;
        RECT 0 36.5 4 39.5 ;
      LAYER METS1 ;
        RECT 0 36.5 4 39.5 ;
      LAYER METS2 ;
        RECT 0 36.5 4 39.5 ;
      LAYER METS3 ;
        RECT 0 36.5 4 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 4 47.5 ;
      LAYER MET6 ;
        RECT 0 44.5 4 47.5 ;
      LAYER METG1 ;
        RECT 0 44.5 4 47.5 ;
      LAYER METS1 ;
        RECT 0 44.5 4 47.5 ;
      LAYER METS2 ;
        RECT 0 44.5 4 47.5 ;
      LAYER METS3 ;
        RECT 0 44.5 4 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 4 55.5 ;
      LAYER MET6 ;
        RECT 0 52.5 4 55.5 ;
      LAYER METG1 ;
        RECT 0 52.5 4 55.5 ;
      LAYER METS1 ;
        RECT 0 52.5 4 55.5 ;
      LAYER METS2 ;
        RECT 0 52.5 4 55.5 ;
      LAYER METS3 ;
        RECT 0 52.5 4 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 4 63.5 ;
      LAYER MET6 ;
        RECT 0 60.5 4 63.5 ;
      LAYER METG1 ;
        RECT 0 60.5 4 63.5 ;
      LAYER METS1 ;
        RECT 0 60.5 4 63.5 ;
      LAYER METS2 ;
        RECT 0 60.5 4 63.5 ;
      LAYER METS3 ;
        RECT 0 60.5 4 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 4 71.5 ;
      LAYER MET6 ;
        RECT 0 68.5 4 71.5 ;
      LAYER METG1 ;
        RECT 0 68.5 4 71.5 ;
      LAYER METS1 ;
        RECT 0 68.5 4 71.5 ;
      LAYER METS2 ;
        RECT 0 68.5 4 71.5 ;
      LAYER METS3 ;
        RECT 0 68.5 4 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 4 103.5 ;
      LAYER MET6 ;
        RECT 0 100.5 4 103.5 ;
      LAYER METG1 ;
        RECT 0 100.5 4 103.5 ;
      LAYER METS1 ;
        RECT 0 100.5 4 103.5 ;
      LAYER METS2 ;
        RECT 0 100.5 4 103.5 ;
      LAYER METS3 ;
        RECT 0 100.5 4 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 4 135.5 ;
      LAYER MET6 ;
        RECT 0 132.5 4 135.5 ;
      LAYER METG1 ;
        RECT 0 132.5 4 135.5 ;
      LAYER METS1 ;
        RECT 0 132.5 4 135.5 ;
      LAYER METS2 ;
        RECT 0 132.5 4 135.5 ;
      LAYER METS3 ;
        RECT 0 132.5 4 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 103.6 4 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 4 107.5 ;
      LAYER MET6 ;
        RECT 0 104.5 4 107.5 ;
      LAYER METG1 ;
        RECT 0 104.5 4 107.5 ;
      LAYER METS1 ;
        RECT 0 104.5 4 107.5 ;
      LAYER METS2 ;
        RECT 0 104.5 4 107.5 ;
      LAYER METS3 ;
        RECT 0 104.5 4 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 4 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 4 115.5 ;
      LAYER MET6 ;
        RECT 0 112.5 4 115.5 ;
      LAYER METG1 ;
        RECT 0 112.5 4 115.5 ;
      LAYER METS1 ;
        RECT 0 112.5 4 115.5 ;
      LAYER METS2 ;
        RECT 0 112.5 4 115.5 ;
      LAYER METS3 ;
        RECT 0 112.5 4 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 4 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 4 119.5 ;
      LAYER MET6 ;
        RECT 0 116.5 4 119.5 ;
      LAYER METG1 ;
        RECT 0 116.5 4 119.5 ;
      LAYER METS1 ;
        RECT 0 116.5 4 119.5 ;
      LAYER METS2 ;
        RECT 0 116.5 4 119.5 ;
      LAYER METS3 ;
        RECT 0 116.5 4 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 4 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 4 123.5 ;
      LAYER MET6 ;
        RECT 0 120.5 4 123.5 ;
      LAYER METG1 ;
        RECT 0 120.5 4 123.5 ;
      LAYER METS1 ;
        RECT 0 120.5 4 123.5 ;
      LAYER METS2 ;
        RECT 0 120.5 4 123.5 ;
      LAYER METS3 ;
        RECT 0 120.5 4 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 4 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 4 127.5 ;
      LAYER MET6 ;
        RECT 0 124.5 4 127.5 ;
      LAYER METG1 ;
        RECT 0 124.5 4 127.5 ;
      LAYER METS1 ;
        RECT 0 124.5 4 127.5 ;
      LAYER METS2 ;
        RECT 0 124.5 4 127.5 ;
      LAYER METS3 ;
        RECT 0 124.5 4 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 4 143.5 ;
      LAYER MET6 ;
        RECT 0 140.5 4 143.5 ;
      LAYER METG1 ;
        RECT 0 140.5 4 143.5 ;
      LAYER METS1 ;
        RECT 0 140.5 4 143.5 ;
      LAYER METS2 ;
        RECT 0 140.5 4 143.5 ;
      LAYER METS3 ;
        RECT 0 140.5 4 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 4 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 4 147.5 ;
      LAYER MET6 ;
        RECT 0 144.5 4 147.5 ;
      LAYER METG1 ;
        RECT 0 144.5 4 147.5 ;
      LAYER METS1 ;
        RECT 0 144.5 4 147.5 ;
      LAYER METS2 ;
        RECT 0 144.5 4 147.5 ;
      LAYER METS3 ;
        RECT 0 144.5 4 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 4 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 4 151.5 ;
      LAYER MET6 ;
        RECT 0 148.5 4 151.5 ;
      LAYER METG1 ;
        RECT 0 148.5 4 151.5 ;
      LAYER METS1 ;
        RECT 0 148.5 4 151.5 ;
      LAYER METS2 ;
        RECT 0 148.5 4 151.5 ;
      LAYER METS3 ;
        RECT 0 148.5 4 151.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 4 110.6 ;
    END
  END VSS
  OBS
    LAYER MET1 ;
      RECT 0 0 4 170 ;
    LAYER CUT12 ;
      RECT 0 0 4 170 ;
    LAYER MET2 ;
      RECT 0 0 4 170 ;
    LAYER CUT23 ;
      RECT 0 0 4 170 ;
    LAYER MET3 ;
      RECT 0 0 4 170 ;
    LAYER CUT34 ;
      RECT 0 0 4 170 ;
    LAYER MET4 ;
      RECT 0 0 4 170 ;
    LAYER CUT45 ;
      RECT 0 0 4 170 ;
    LAYER MET5 ;
      RECT 0 0 4 170 ;
    LAYER CUT56 ;
      RECT 0 0 4 170 ;
    LAYER MET6 ;
      RECT 0 0 4 170 ;
    LAYER CUTS1 ;
      RECT 0 0 4 170 ;
    LAYER METS1 ;
      RECT 0 0 4 170 ;
    LAYER CUTS2 ;
      RECT 0 0 4 170 ;
    LAYER METS2 ;
      RECT 0 0 4 170 ;
    LAYER CUTS3 ;
      RECT 0 0 4 170 ;
    LAYER METS3 ;
      RECT 0 0 4 170 ;
    LAYER CUTG1 ;
      RECT 0 0 4 170 ;
    LAYER METG1 ;
      RECT 0 0 4 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 4.000 2.000 ;
  END
END IOCB2EDC2E4C01


MACRO IOCB2ES14C0A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2ES14C0A1 0 0 ;
  SIZE 1 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 28.5 1 31.5 ;
      LAYER MET6 ;
        RECT 0 28.5 1 31.5 ;
      LAYER METG1 ;
        RECT 0 28.5 1 31.5 ;
      LAYER METS1 ;
        RECT 0 28.5 1 31.5 ;
      LAYER METS2 ;
        RECT 0 28.5 1 31.5 ;
      LAYER METS3 ;
        RECT 0 28.5 1 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 1 35.5 ;
      LAYER MET6 ;
        RECT 0 32.5 1 35.5 ;
      LAYER METG1 ;
        RECT 0 32.5 1 35.5 ;
      LAYER METS1 ;
        RECT 0 32.5 1 35.5 ;
      LAYER METS2 ;
        RECT 0 32.5 1 35.5 ;
      LAYER METS3 ;
        RECT 0 32.5 1 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 1 43.5 ;
      LAYER MET6 ;
        RECT 0 40.5 1 43.5 ;
      LAYER METG1 ;
        RECT 0 40.5 1 43.5 ;
      LAYER METS1 ;
        RECT 0 40.5 1 43.5 ;
      LAYER METS2 ;
        RECT 0 40.5 1 43.5 ;
      LAYER METS3 ;
        RECT 0 40.5 1 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 1 51.5 ;
      LAYER MET6 ;
        RECT 0 48.5 1 51.5 ;
      LAYER METG1 ;
        RECT 0 48.5 1 51.5 ;
      LAYER METS1 ;
        RECT 0 48.5 1 51.5 ;
      LAYER METS2 ;
        RECT 0 48.5 1 51.5 ;
      LAYER METS3 ;
        RECT 0 48.5 1 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 1 59.5 ;
      LAYER MET6 ;
        RECT 0 56.5 1 59.5 ;
      LAYER METG1 ;
        RECT 0 56.5 1 59.5 ;
      LAYER METS1 ;
        RECT 0 56.5 1 59.5 ;
      LAYER METS2 ;
        RECT 0 56.5 1 59.5 ;
      LAYER METS3 ;
        RECT 0 56.5 1 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 1 67.5 ;
      LAYER MET6 ;
        RECT 0 64.5 1 67.5 ;
      LAYER METG1 ;
        RECT 0 64.5 1 67.5 ;
      LAYER METS1 ;
        RECT 0 64.5 1 67.5 ;
      LAYER METS2 ;
        RECT 0 64.5 1 67.5 ;
      LAYER METS3 ;
        RECT 0 64.5 1 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 1 75.5 ;
      LAYER MET6 ;
        RECT 0 72.5 1 75.5 ;
      LAYER METG1 ;
        RECT 0 72.5 1 75.5 ;
      LAYER METS1 ;
        RECT 0 72.5 1 75.5 ;
      LAYER METS2 ;
        RECT 0 72.5 1 75.5 ;
      LAYER METS3 ;
        RECT 0 72.5 1 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 1 111.5 ;
      LAYER MET6 ;
        RECT 0 108.5 1 111.5 ;
      LAYER METG1 ;
        RECT 0 108.5 1 111.5 ;
      LAYER METS1 ;
        RECT 0 108.5 1 111.5 ;
      LAYER METS2 ;
        RECT 0 108.5 1 111.5 ;
      LAYER METS3 ;
        RECT 0 108.5 1 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 1 131.5 ;
      LAYER MET6 ;
        RECT 0 128.5 1 131.5 ;
      LAYER METG1 ;
        RECT 0 128.5 1 131.5 ;
      LAYER METS1 ;
        RECT 0 128.5 1 131.5 ;
      LAYER METS2 ;
        RECT 0 128.5 1 131.5 ;
      LAYER METS3 ;
        RECT 0 128.5 1 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 1 139.5 ;
      LAYER MET6 ;
        RECT 0 136.5 1 139.5 ;
      LAYER METG1 ;
        RECT 0 136.5 1 139.5 ;
      LAYER METS1 ;
        RECT 0 136.5 1 139.5 ;
      LAYER METS2 ;
        RECT 0 136.5 1 139.5 ;
      LAYER METS3 ;
        RECT 0 136.5 1 139.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 75.6 1 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 1 79.5 ;
      LAYER MET6 ;
        RECT 0 76.5 1 79.5 ;
      LAYER METG1 ;
        RECT 0 76.5 1 79.5 ;
      LAYER METS1 ;
        RECT 0 76.5 1 79.5 ;
      LAYER METS2 ;
        RECT 0 76.5 1 79.5 ;
      LAYER METS3 ;
        RECT 0 76.5 1 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 1 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 1 83.5 ;
      LAYER MET6 ;
        RECT 0 80.5 1 83.5 ;
      LAYER METG1 ;
        RECT 0 80.5 1 83.5 ;
      LAYER METS1 ;
        RECT 0 80.5 1 83.5 ;
      LAYER METS2 ;
        RECT 0 80.5 1 83.5 ;
      LAYER METS3 ;
        RECT 0 80.5 1 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 1 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 1 87.5 ;
      LAYER MET6 ;
        RECT 0 84.5 1 87.5 ;
      LAYER METG1 ;
        RECT 0 84.5 1 87.5 ;
      LAYER METS1 ;
        RECT 0 84.5 1 87.5 ;
      LAYER METS2 ;
        RECT 0 84.5 1 87.5 ;
      LAYER METS3 ;
        RECT 0 84.5 1 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 1 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 1 91.5 ;
      LAYER MET6 ;
        RECT 0 88.5 1 91.5 ;
      LAYER METG1 ;
        RECT 0 88.5 1 91.5 ;
      LAYER METS1 ;
        RECT 0 88.5 1 91.5 ;
      LAYER METS2 ;
        RECT 0 88.5 1 91.5 ;
      LAYER METS3 ;
        RECT 0 88.5 1 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 1 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 1 95.5 ;
      LAYER MET6 ;
        RECT 0 92.5 1 95.5 ;
      LAYER METG1 ;
        RECT 0 92.5 1 95.5 ;
      LAYER METS1 ;
        RECT 0 92.5 1 95.5 ;
      LAYER METS2 ;
        RECT 0 92.5 1 95.5 ;
      LAYER METS3 ;
        RECT 0 92.5 1 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 1 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 1 99.5 ;
      LAYER MET6 ;
        RECT 0 96.5 1 99.5 ;
      LAYER METG1 ;
        RECT 0 96.5 1 99.5 ;
      LAYER METS1 ;
        RECT 0 96.5 1 99.5 ;
      LAYER METS2 ;
        RECT 0 96.5 1 99.5 ;
      LAYER METS3 ;
        RECT 0 96.5 1 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 1 155.5 ;
      LAYER MET6 ;
        RECT 0 152.5 1 155.5 ;
      LAYER METG1 ;
        RECT 0 152.5 1 155.5 ;
      LAYER METS1 ;
        RECT 0 152.5 1 155.5 ;
      LAYER METS2 ;
        RECT 0 152.5 1 155.5 ;
      LAYER METS3 ;
        RECT 0 152.5 1 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 1 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 1 159.5 ;
      LAYER MET6 ;
        RECT 0 156.5 1 159.5 ;
      LAYER METG1 ;
        RECT 0 156.5 1 159.5 ;
      LAYER METS1 ;
        RECT 0 156.5 1 159.5 ;
      LAYER METS2 ;
        RECT 0 156.5 1 159.5 ;
      LAYER METS3 ;
        RECT 0 156.5 1 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 1 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 1 163.5 ;
      LAYER MET6 ;
        RECT 0 160.5 1 163.5 ;
      LAYER METG1 ;
        RECT 0 160.5 1 163.5 ;
      LAYER METS1 ;
        RECT 0 160.5 1 163.5 ;
      LAYER METS2 ;
        RECT 0 160.5 1 163.5 ;
      LAYER METS3 ;
        RECT 0 160.5 1 163.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 4.5 1 7.5 ;
      LAYER MET6 ;
        RECT 0 4.5 1 7.5 ;
      LAYER METG1 ;
        RECT 0 4.5 1 7.5 ;
      LAYER METS1 ;
        RECT 0 4.5 1 7.5 ;
      LAYER METS2 ;
        RECT 0 4.5 1 7.5 ;
      LAYER METS3 ;
        RECT 0 4.5 1 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 1 11.5 ;
      LAYER MET6 ;
        RECT 0 8.5 1 11.5 ;
      LAYER METG1 ;
        RECT 0 8.5 1 11.5 ;
      LAYER METS1 ;
        RECT 0 8.5 1 11.5 ;
      LAYER METS2 ;
        RECT 0 8.5 1 11.5 ;
      LAYER METS3 ;
        RECT 0 8.5 1 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 1 23.5 ;
      LAYER MET6 ;
        RECT 0 20.5 1 23.5 ;
      LAYER METG1 ;
        RECT 0 20.5 1 23.5 ;
      LAYER METS1 ;
        RECT 0 20.5 1 23.5 ;
      LAYER METS2 ;
        RECT 0 20.5 1 23.5 ;
      LAYER METS3 ;
        RECT 0 20.5 1 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 1 27.5 ;
      LAYER MET6 ;
        RECT 0 24.5 1 27.5 ;
      LAYER METG1 ;
        RECT 0 24.5 1 27.5 ;
      LAYER METS1 ;
        RECT 0 24.5 1 27.5 ;
      LAYER METS2 ;
        RECT 0 24.5 1 27.5 ;
      LAYER METS3 ;
        RECT 0 24.5 1 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 1 39.5 ;
      LAYER MET6 ;
        RECT 0 36.5 1 39.5 ;
      LAYER METG1 ;
        RECT 0 36.5 1 39.5 ;
      LAYER METS1 ;
        RECT 0 36.5 1 39.5 ;
      LAYER METS2 ;
        RECT 0 36.5 1 39.5 ;
      LAYER METS3 ;
        RECT 0 36.5 1 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 1 47.5 ;
      LAYER MET6 ;
        RECT 0 44.5 1 47.5 ;
      LAYER METG1 ;
        RECT 0 44.5 1 47.5 ;
      LAYER METS1 ;
        RECT 0 44.5 1 47.5 ;
      LAYER METS2 ;
        RECT 0 44.5 1 47.5 ;
      LAYER METS3 ;
        RECT 0 44.5 1 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 1 55.5 ;
      LAYER MET6 ;
        RECT 0 52.5 1 55.5 ;
      LAYER METG1 ;
        RECT 0 52.5 1 55.5 ;
      LAYER METS1 ;
        RECT 0 52.5 1 55.5 ;
      LAYER METS2 ;
        RECT 0 52.5 1 55.5 ;
      LAYER METS3 ;
        RECT 0 52.5 1 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 1 63.5 ;
      LAYER MET6 ;
        RECT 0 60.5 1 63.5 ;
      LAYER METG1 ;
        RECT 0 60.5 1 63.5 ;
      LAYER METS1 ;
        RECT 0 60.5 1 63.5 ;
      LAYER METS2 ;
        RECT 0 60.5 1 63.5 ;
      LAYER METS3 ;
        RECT 0 60.5 1 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 1 71.5 ;
      LAYER MET6 ;
        RECT 0 68.5 1 71.5 ;
      LAYER METG1 ;
        RECT 0 68.5 1 71.5 ;
      LAYER METS1 ;
        RECT 0 68.5 1 71.5 ;
      LAYER METS2 ;
        RECT 0 68.5 1 71.5 ;
      LAYER METS3 ;
        RECT 0 68.5 1 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 1 103.5 ;
      LAYER MET6 ;
        RECT 0 100.5 1 103.5 ;
      LAYER METG1 ;
        RECT 0 100.5 1 103.5 ;
      LAYER METS1 ;
        RECT 0 100.5 1 103.5 ;
      LAYER METS2 ;
        RECT 0 100.5 1 103.5 ;
      LAYER METS3 ;
        RECT 0 100.5 1 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 1 135.5 ;
      LAYER MET6 ;
        RECT 0 132.5 1 135.5 ;
      LAYER METG1 ;
        RECT 0 132.5 1 135.5 ;
      LAYER METS1 ;
        RECT 0 132.5 1 135.5 ;
      LAYER METS2 ;
        RECT 0 132.5 1 135.5 ;
      LAYER METS3 ;
        RECT 0 132.5 1 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 103.6 1 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 1 107.5 ;
      LAYER MET6 ;
        RECT 0 104.5 1 107.5 ;
      LAYER METG1 ;
        RECT 0 104.5 1 107.5 ;
      LAYER METS1 ;
        RECT 0 104.5 1 107.5 ;
      LAYER METS2 ;
        RECT 0 104.5 1 107.5 ;
      LAYER METS3 ;
        RECT 0 104.5 1 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 1 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 1 115.5 ;
      LAYER MET6 ;
        RECT 0 112.5 1 115.5 ;
      LAYER METG1 ;
        RECT 0 112.5 1 115.5 ;
      LAYER METS1 ;
        RECT 0 112.5 1 115.5 ;
      LAYER METS2 ;
        RECT 0 112.5 1 115.5 ;
      LAYER METS3 ;
        RECT 0 112.5 1 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 1 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 1 119.5 ;
      LAYER MET6 ;
        RECT 0 116.5 1 119.5 ;
      LAYER METG1 ;
        RECT 0 116.5 1 119.5 ;
      LAYER METS1 ;
        RECT 0 116.5 1 119.5 ;
      LAYER METS2 ;
        RECT 0 116.5 1 119.5 ;
      LAYER METS3 ;
        RECT 0 116.5 1 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 1 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 1 123.5 ;
      LAYER MET6 ;
        RECT 0 120.5 1 123.5 ;
      LAYER METG1 ;
        RECT 0 120.5 1 123.5 ;
      LAYER METS1 ;
        RECT 0 120.5 1 123.5 ;
      LAYER METS2 ;
        RECT 0 120.5 1 123.5 ;
      LAYER METS3 ;
        RECT 0 120.5 1 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 1 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 1 127.5 ;
      LAYER MET6 ;
        RECT 0 124.5 1 127.5 ;
      LAYER METG1 ;
        RECT 0 124.5 1 127.5 ;
      LAYER METS1 ;
        RECT 0 124.5 1 127.5 ;
      LAYER METS2 ;
        RECT 0 124.5 1 127.5 ;
      LAYER METS3 ;
        RECT 0 124.5 1 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 1 143.5 ;
      LAYER MET6 ;
        RECT 0 140.5 1 143.5 ;
      LAYER METG1 ;
        RECT 0 140.5 1 143.5 ;
      LAYER METS1 ;
        RECT 0 140.5 1 143.5 ;
      LAYER METS2 ;
        RECT 0 140.5 1 143.5 ;
      LAYER METS3 ;
        RECT 0 140.5 1 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 1 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 1 147.5 ;
      LAYER MET6 ;
        RECT 0 144.5 1 147.5 ;
      LAYER METG1 ;
        RECT 0 144.5 1 147.5 ;
      LAYER METS1 ;
        RECT 0 144.5 1 147.5 ;
      LAYER METS2 ;
        RECT 0 144.5 1 147.5 ;
      LAYER METS3 ;
        RECT 0 144.5 1 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 1 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 1 151.5 ;
      LAYER MET6 ;
        RECT 0 148.5 1 151.5 ;
      LAYER METG1 ;
        RECT 0 148.5 1 151.5 ;
      LAYER METS1 ;
        RECT 0 148.5 1 151.5 ;
      LAYER METS2 ;
        RECT 0 148.5 1 151.5 ;
      LAYER METS3 ;
        RECT 0 148.5 1 151.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 1 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 1 15.5 ;
      LAYER MET6 ;
        RECT 0 12.5 1 15.5 ;
      LAYER METG1 ;
        RECT 0 12.5 1 15.5 ;
      LAYER METS1 ;
        RECT 0 12.5 1 15.5 ;
      LAYER METS2 ;
        RECT 0 12.5 1 15.5 ;
      LAYER METS3 ;
        RECT 0 12.5 1 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 1 19.5 ;
      LAYER MET6 ;
        RECT 0 16.5 1 19.5 ;
      LAYER METG1 ;
        RECT 0 16.5 1 19.5 ;
      LAYER METS1 ;
        RECT 0 16.5 1 19.5 ;
      LAYER METS2 ;
        RECT 0 16.5 1 19.5 ;
      LAYER METS3 ;
        RECT 0 16.5 1 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 1 170 ;
    LAYER CUT12 ;
      RECT 0 0 1 170 ;
    LAYER MET2 ;
      RECT 0 0 1 170 ;
    LAYER CUT23 ;
      RECT 0 0 1 170 ;
    LAYER MET3 ;
      RECT 0 0 1 170 ;
    LAYER CUT34 ;
      RECT 0 0 1 170 ;
    LAYER MET4 ;
      RECT 0 0 1 170 ;
    LAYER CUT45 ;
      RECT 0 0 1 170 ;
    LAYER MET5 ;
      RECT 0 0 1 170 ;
    LAYER CUT56 ;
      RECT 0 0 1 170 ;
    LAYER MET6 ;
      RECT 0 0 1 170 ;
    LAYER CUTS1 ;
      RECT 0 0 1 170 ;
    LAYER METS1 ;
      RECT 0 0 1 170 ;
    LAYER CUTS2 ;
      RECT 0 0 1 170 ;
    LAYER METS2 ;
      RECT 0 0 1 170 ;
    LAYER CUTS3 ;
      RECT 0 0 1 170 ;
    LAYER METS3 ;
      RECT 0 0 1 170 ;
    LAYER CUTG1 ;
      RECT 0 0 1 170 ;
    LAYER METG1 ;
      RECT 0 0 1 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 1.000 2.000 ;
  END
END IOCB2ES14C0A1


MACRO IOCB2ES24C0A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2ES24C0A1 0 0 ;
  SIZE 2 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 28.5 2 31.5 ;
      LAYER MET6 ;
        RECT 0 28.5 2 31.5 ;
      LAYER METG1 ;
        RECT 0 28.5 2 31.5 ;
      LAYER METS1 ;
        RECT 0 28.5 2 31.5 ;
      LAYER METS2 ;
        RECT 0 28.5 2 31.5 ;
      LAYER METS3 ;
        RECT 0 28.5 2 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 2 35.5 ;
      LAYER MET6 ;
        RECT 0 32.5 2 35.5 ;
      LAYER METG1 ;
        RECT 0 32.5 2 35.5 ;
      LAYER METS1 ;
        RECT 0 32.5 2 35.5 ;
      LAYER METS2 ;
        RECT 0 32.5 2 35.5 ;
      LAYER METS3 ;
        RECT 0 32.5 2 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 2 43.5 ;
      LAYER MET6 ;
        RECT 0 40.5 2 43.5 ;
      LAYER METG1 ;
        RECT 0 40.5 2 43.5 ;
      LAYER METS1 ;
        RECT 0 40.5 2 43.5 ;
      LAYER METS2 ;
        RECT 0 40.5 2 43.5 ;
      LAYER METS3 ;
        RECT 0 40.5 2 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 2 51.5 ;
      LAYER MET6 ;
        RECT 0 48.5 2 51.5 ;
      LAYER METG1 ;
        RECT 0 48.5 2 51.5 ;
      LAYER METS1 ;
        RECT 0 48.5 2 51.5 ;
      LAYER METS2 ;
        RECT 0 48.5 2 51.5 ;
      LAYER METS3 ;
        RECT 0 48.5 2 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 2 59.5 ;
      LAYER MET6 ;
        RECT 0 56.5 2 59.5 ;
      LAYER METG1 ;
        RECT 0 56.5 2 59.5 ;
      LAYER METS1 ;
        RECT 0 56.5 2 59.5 ;
      LAYER METS2 ;
        RECT 0 56.5 2 59.5 ;
      LAYER METS3 ;
        RECT 0 56.5 2 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 2 67.5 ;
      LAYER MET6 ;
        RECT 0 64.5 2 67.5 ;
      LAYER METG1 ;
        RECT 0 64.5 2 67.5 ;
      LAYER METS1 ;
        RECT 0 64.5 2 67.5 ;
      LAYER METS2 ;
        RECT 0 64.5 2 67.5 ;
      LAYER METS3 ;
        RECT 0 64.5 2 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 2 75.5 ;
      LAYER MET6 ;
        RECT 0 72.5 2 75.5 ;
      LAYER METG1 ;
        RECT 0 72.5 2 75.5 ;
      LAYER METS1 ;
        RECT 0 72.5 2 75.5 ;
      LAYER METS2 ;
        RECT 0 72.5 2 75.5 ;
      LAYER METS3 ;
        RECT 0 72.5 2 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 2 111.5 ;
      LAYER MET6 ;
        RECT 0 108.5 2 111.5 ;
      LAYER METG1 ;
        RECT 0 108.5 2 111.5 ;
      LAYER METS1 ;
        RECT 0 108.5 2 111.5 ;
      LAYER METS2 ;
        RECT 0 108.5 2 111.5 ;
      LAYER METS3 ;
        RECT 0 108.5 2 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 2 131.5 ;
      LAYER MET6 ;
        RECT 0 128.5 2 131.5 ;
      LAYER METG1 ;
        RECT 0 128.5 2 131.5 ;
      LAYER METS1 ;
        RECT 0 128.5 2 131.5 ;
      LAYER METS2 ;
        RECT 0 128.5 2 131.5 ;
      LAYER METS3 ;
        RECT 0 128.5 2 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 2 139.5 ;
      LAYER MET6 ;
        RECT 0 136.5 2 139.5 ;
      LAYER METG1 ;
        RECT 0 136.5 2 139.5 ;
      LAYER METS1 ;
        RECT 0 136.5 2 139.5 ;
      LAYER METS2 ;
        RECT 0 136.5 2 139.5 ;
      LAYER METS3 ;
        RECT 0 136.5 2 139.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 75.6 2 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 2 79.5 ;
      LAYER MET6 ;
        RECT 0 76.5 2 79.5 ;
      LAYER METG1 ;
        RECT 0 76.5 2 79.5 ;
      LAYER METS1 ;
        RECT 0 76.5 2 79.5 ;
      LAYER METS2 ;
        RECT 0 76.5 2 79.5 ;
      LAYER METS3 ;
        RECT 0 76.5 2 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 2 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 2 83.5 ;
      LAYER MET6 ;
        RECT 0 80.5 2 83.5 ;
      LAYER METG1 ;
        RECT 0 80.5 2 83.5 ;
      LAYER METS1 ;
        RECT 0 80.5 2 83.5 ;
      LAYER METS2 ;
        RECT 0 80.5 2 83.5 ;
      LAYER METS3 ;
        RECT 0 80.5 2 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 2 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 2 87.5 ;
      LAYER MET6 ;
        RECT 0 84.5 2 87.5 ;
      LAYER METG1 ;
        RECT 0 84.5 2 87.5 ;
      LAYER METS1 ;
        RECT 0 84.5 2 87.5 ;
      LAYER METS2 ;
        RECT 0 84.5 2 87.5 ;
      LAYER METS3 ;
        RECT 0 84.5 2 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 2 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 2 91.5 ;
      LAYER MET6 ;
        RECT 0 88.5 2 91.5 ;
      LAYER METG1 ;
        RECT 0 88.5 2 91.5 ;
      LAYER METS1 ;
        RECT 0 88.5 2 91.5 ;
      LAYER METS2 ;
        RECT 0 88.5 2 91.5 ;
      LAYER METS3 ;
        RECT 0 88.5 2 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 2 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 2 95.5 ;
      LAYER MET6 ;
        RECT 0 92.5 2 95.5 ;
      LAYER METG1 ;
        RECT 0 92.5 2 95.5 ;
      LAYER METS1 ;
        RECT 0 92.5 2 95.5 ;
      LAYER METS2 ;
        RECT 0 92.5 2 95.5 ;
      LAYER METS3 ;
        RECT 0 92.5 2 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 2 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 2 99.5 ;
      LAYER MET6 ;
        RECT 0 96.5 2 99.5 ;
      LAYER METG1 ;
        RECT 0 96.5 2 99.5 ;
      LAYER METS1 ;
        RECT 0 96.5 2 99.5 ;
      LAYER METS2 ;
        RECT 0 96.5 2 99.5 ;
      LAYER METS3 ;
        RECT 0 96.5 2 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 2 155.5 ;
      LAYER MET6 ;
        RECT 0 152.5 2 155.5 ;
      LAYER METG1 ;
        RECT 0 152.5 2 155.5 ;
      LAYER METS1 ;
        RECT 0 152.5 2 155.5 ;
      LAYER METS2 ;
        RECT 0 152.5 2 155.5 ;
      LAYER METS3 ;
        RECT 0 152.5 2 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 2 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 2 159.5 ;
      LAYER MET6 ;
        RECT 0 156.5 2 159.5 ;
      LAYER METG1 ;
        RECT 0 156.5 2 159.5 ;
      LAYER METS1 ;
        RECT 0 156.5 2 159.5 ;
      LAYER METS2 ;
        RECT 0 156.5 2 159.5 ;
      LAYER METS3 ;
        RECT 0 156.5 2 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 2 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 2 163.5 ;
      LAYER MET6 ;
        RECT 0 160.5 2 163.5 ;
      LAYER METG1 ;
        RECT 0 160.5 2 163.5 ;
      LAYER METS1 ;
        RECT 0 160.5 2 163.5 ;
      LAYER METS2 ;
        RECT 0 160.5 2 163.5 ;
      LAYER METS3 ;
        RECT 0 160.5 2 163.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 4.5 2 7.5 ;
      LAYER MET6 ;
        RECT 0 4.5 2 7.5 ;
      LAYER METG1 ;
        RECT 0 4.5 2 7.5 ;
      LAYER METS1 ;
        RECT 0 4.5 2 7.5 ;
      LAYER METS2 ;
        RECT 0 4.5 2 7.5 ;
      LAYER METS3 ;
        RECT 0 4.5 2 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 2 11.5 ;
      LAYER MET6 ;
        RECT 0 8.5 2 11.5 ;
      LAYER METG1 ;
        RECT 0 8.5 2 11.5 ;
      LAYER METS1 ;
        RECT 0 8.5 2 11.5 ;
      LAYER METS2 ;
        RECT 0 8.5 2 11.5 ;
      LAYER METS3 ;
        RECT 0 8.5 2 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 2 23.5 ;
      LAYER MET6 ;
        RECT 0 20.5 2 23.5 ;
      LAYER METG1 ;
        RECT 0 20.5 2 23.5 ;
      LAYER METS1 ;
        RECT 0 20.5 2 23.5 ;
      LAYER METS2 ;
        RECT 0 20.5 2 23.5 ;
      LAYER METS3 ;
        RECT 0 20.5 2 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 2 27.5 ;
      LAYER MET6 ;
        RECT 0 24.5 2 27.5 ;
      LAYER METG1 ;
        RECT 0 24.5 2 27.5 ;
      LAYER METS1 ;
        RECT 0 24.5 2 27.5 ;
      LAYER METS2 ;
        RECT 0 24.5 2 27.5 ;
      LAYER METS3 ;
        RECT 0 24.5 2 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 2 39.5 ;
      LAYER MET6 ;
        RECT 0 36.5 2 39.5 ;
      LAYER METG1 ;
        RECT 0 36.5 2 39.5 ;
      LAYER METS1 ;
        RECT 0 36.5 2 39.5 ;
      LAYER METS2 ;
        RECT 0 36.5 2 39.5 ;
      LAYER METS3 ;
        RECT 0 36.5 2 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 2 47.5 ;
      LAYER MET6 ;
        RECT 0 44.5 2 47.5 ;
      LAYER METG1 ;
        RECT 0 44.5 2 47.5 ;
      LAYER METS1 ;
        RECT 0 44.5 2 47.5 ;
      LAYER METS2 ;
        RECT 0 44.5 2 47.5 ;
      LAYER METS3 ;
        RECT 0 44.5 2 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 2 55.5 ;
      LAYER MET6 ;
        RECT 0 52.5 2 55.5 ;
      LAYER METG1 ;
        RECT 0 52.5 2 55.5 ;
      LAYER METS1 ;
        RECT 0 52.5 2 55.5 ;
      LAYER METS2 ;
        RECT 0 52.5 2 55.5 ;
      LAYER METS3 ;
        RECT 0 52.5 2 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 2 63.5 ;
      LAYER MET6 ;
        RECT 0 60.5 2 63.5 ;
      LAYER METG1 ;
        RECT 0 60.5 2 63.5 ;
      LAYER METS1 ;
        RECT 0 60.5 2 63.5 ;
      LAYER METS2 ;
        RECT 0 60.5 2 63.5 ;
      LAYER METS3 ;
        RECT 0 60.5 2 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 2 71.5 ;
      LAYER MET6 ;
        RECT 0 68.5 2 71.5 ;
      LAYER METG1 ;
        RECT 0 68.5 2 71.5 ;
      LAYER METS1 ;
        RECT 0 68.5 2 71.5 ;
      LAYER METS2 ;
        RECT 0 68.5 2 71.5 ;
      LAYER METS3 ;
        RECT 0 68.5 2 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 2 103.5 ;
      LAYER MET6 ;
        RECT 0 100.5 2 103.5 ;
      LAYER METG1 ;
        RECT 0 100.5 2 103.5 ;
      LAYER METS1 ;
        RECT 0 100.5 2 103.5 ;
      LAYER METS2 ;
        RECT 0 100.5 2 103.5 ;
      LAYER METS3 ;
        RECT 0 100.5 2 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 2 135.5 ;
      LAYER MET6 ;
        RECT 0 132.5 2 135.5 ;
      LAYER METG1 ;
        RECT 0 132.5 2 135.5 ;
      LAYER METS1 ;
        RECT 0 132.5 2 135.5 ;
      LAYER METS2 ;
        RECT 0 132.5 2 135.5 ;
      LAYER METS3 ;
        RECT 0 132.5 2 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 103.6 2 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 2 107.5 ;
      LAYER MET6 ;
        RECT 0 104.5 2 107.5 ;
      LAYER METG1 ;
        RECT 0 104.5 2 107.5 ;
      LAYER METS1 ;
        RECT 0 104.5 2 107.5 ;
      LAYER METS2 ;
        RECT 0 104.5 2 107.5 ;
      LAYER METS3 ;
        RECT 0 104.5 2 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 2 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 2 115.5 ;
      LAYER MET6 ;
        RECT 0 112.5 2 115.5 ;
      LAYER METG1 ;
        RECT 0 112.5 2 115.5 ;
      LAYER METS1 ;
        RECT 0 112.5 2 115.5 ;
      LAYER METS2 ;
        RECT 0 112.5 2 115.5 ;
      LAYER METS3 ;
        RECT 0 112.5 2 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 2 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 2 119.5 ;
      LAYER MET6 ;
        RECT 0 116.5 2 119.5 ;
      LAYER METG1 ;
        RECT 0 116.5 2 119.5 ;
      LAYER METS1 ;
        RECT 0 116.5 2 119.5 ;
      LAYER METS2 ;
        RECT 0 116.5 2 119.5 ;
      LAYER METS3 ;
        RECT 0 116.5 2 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 2 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 2 123.5 ;
      LAYER MET6 ;
        RECT 0 120.5 2 123.5 ;
      LAYER METG1 ;
        RECT 0 120.5 2 123.5 ;
      LAYER METS1 ;
        RECT 0 120.5 2 123.5 ;
      LAYER METS2 ;
        RECT 0 120.5 2 123.5 ;
      LAYER METS3 ;
        RECT 0 120.5 2 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 2 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 2 127.5 ;
      LAYER MET6 ;
        RECT 0 124.5 2 127.5 ;
      LAYER METG1 ;
        RECT 0 124.5 2 127.5 ;
      LAYER METS1 ;
        RECT 0 124.5 2 127.5 ;
      LAYER METS2 ;
        RECT 0 124.5 2 127.5 ;
      LAYER METS3 ;
        RECT 0 124.5 2 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 2 143.5 ;
      LAYER MET6 ;
        RECT 0 140.5 2 143.5 ;
      LAYER METG1 ;
        RECT 0 140.5 2 143.5 ;
      LAYER METS1 ;
        RECT 0 140.5 2 143.5 ;
      LAYER METS2 ;
        RECT 0 140.5 2 143.5 ;
      LAYER METS3 ;
        RECT 0 140.5 2 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 2 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 2 147.5 ;
      LAYER MET6 ;
        RECT 0 144.5 2 147.5 ;
      LAYER METG1 ;
        RECT 0 144.5 2 147.5 ;
      LAYER METS1 ;
        RECT 0 144.5 2 147.5 ;
      LAYER METS2 ;
        RECT 0 144.5 2 147.5 ;
      LAYER METS3 ;
        RECT 0 144.5 2 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 2 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 2 151.5 ;
      LAYER MET6 ;
        RECT 0 148.5 2 151.5 ;
      LAYER METG1 ;
        RECT 0 148.5 2 151.5 ;
      LAYER METS1 ;
        RECT 0 148.5 2 151.5 ;
      LAYER METS2 ;
        RECT 0 148.5 2 151.5 ;
      LAYER METS3 ;
        RECT 0 148.5 2 151.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 2 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 2 15.5 ;
      LAYER MET6 ;
        RECT 0 12.5 2 15.5 ;
      LAYER METG1 ;
        RECT 0 12.5 2 15.5 ;
      LAYER METS1 ;
        RECT 0 12.5 2 15.5 ;
      LAYER METS2 ;
        RECT 0 12.5 2 15.5 ;
      LAYER METS3 ;
        RECT 0 12.5 2 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 2 19.5 ;
      LAYER MET6 ;
        RECT 0 16.5 2 19.5 ;
      LAYER METG1 ;
        RECT 0 16.5 2 19.5 ;
      LAYER METS1 ;
        RECT 0 16.5 2 19.5 ;
      LAYER METS2 ;
        RECT 0 16.5 2 19.5 ;
      LAYER METS3 ;
        RECT 0 16.5 2 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 2 170 ;
    LAYER CUT12 ;
      RECT 0 0 2 170 ;
    LAYER MET2 ;
      RECT 0 0 2 170 ;
    LAYER CUT23 ;
      RECT 0 0 2 170 ;
    LAYER MET3 ;
      RECT 0 0 2 170 ;
    LAYER CUT34 ;
      RECT 0 0 2 170 ;
    LAYER MET4 ;
      RECT 0 0 2 170 ;
    LAYER CUT45 ;
      RECT 0 0 2 170 ;
    LAYER MET5 ;
      RECT 0 0 2 170 ;
    LAYER CUT56 ;
      RECT 0 0 2 170 ;
    LAYER MET6 ;
      RECT 0 0 2 170 ;
    LAYER CUTS1 ;
      RECT 0 0 2 170 ;
    LAYER METS1 ;
      RECT 0 0 2 170 ;
    LAYER CUTS2 ;
      RECT 0 0 2 170 ;
    LAYER METS2 ;
      RECT 0 0 2 170 ;
    LAYER CUTS3 ;
      RECT 0 0 2 170 ;
    LAYER METS3 ;
      RECT 0 0 2 170 ;
    LAYER CUTG1 ;
      RECT 0 0 2 170 ;
    LAYER METG1 ;
      RECT 0 0 2 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 2.000 2.000 ;
  END
END IOCB2ES24C0A1


MACRO IOCB2ES54C0A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2ES54C0A1 0 0 ;
  SIZE 5 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 28.5 5 31.5 ;
      LAYER MET6 ;
        RECT 0 28.5 5 31.5 ;
      LAYER METG1 ;
        RECT 0 28.5 5 31.5 ;
      LAYER METS1 ;
        RECT 0 28.5 5 31.5 ;
      LAYER METS2 ;
        RECT 0 28.5 5 31.5 ;
      LAYER METS3 ;
        RECT 0 28.5 5 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 5 35.5 ;
      LAYER MET6 ;
        RECT 0 32.5 5 35.5 ;
      LAYER METG1 ;
        RECT 0 32.5 5 35.5 ;
      LAYER METS1 ;
        RECT 0 32.5 5 35.5 ;
      LAYER METS2 ;
        RECT 0 32.5 5 35.5 ;
      LAYER METS3 ;
        RECT 0 32.5 5 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 5 43.5 ;
      LAYER MET6 ;
        RECT 0 40.5 5 43.5 ;
      LAYER METG1 ;
        RECT 0 40.5 5 43.5 ;
      LAYER METS1 ;
        RECT 0 40.5 5 43.5 ;
      LAYER METS2 ;
        RECT 0 40.5 5 43.5 ;
      LAYER METS3 ;
        RECT 0 40.5 5 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 5 51.5 ;
      LAYER MET6 ;
        RECT 0 48.5 5 51.5 ;
      LAYER METG1 ;
        RECT 0 48.5 5 51.5 ;
      LAYER METS1 ;
        RECT 0 48.5 5 51.5 ;
      LAYER METS2 ;
        RECT 0 48.5 5 51.5 ;
      LAYER METS3 ;
        RECT 0 48.5 5 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 5 59.5 ;
      LAYER MET6 ;
        RECT 0 56.5 5 59.5 ;
      LAYER METG1 ;
        RECT 0 56.5 5 59.5 ;
      LAYER METS1 ;
        RECT 0 56.5 5 59.5 ;
      LAYER METS2 ;
        RECT 0 56.5 5 59.5 ;
      LAYER METS3 ;
        RECT 0 56.5 5 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 5 67.5 ;
      LAYER MET6 ;
        RECT 0 64.5 5 67.5 ;
      LAYER METG1 ;
        RECT 0 64.5 5 67.5 ;
      LAYER METS1 ;
        RECT 0 64.5 5 67.5 ;
      LAYER METS2 ;
        RECT 0 64.5 5 67.5 ;
      LAYER METS3 ;
        RECT 0 64.5 5 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 5 75.5 ;
      LAYER MET6 ;
        RECT 0 72.5 5 75.5 ;
      LAYER METG1 ;
        RECT 0 72.5 5 75.5 ;
      LAYER METS1 ;
        RECT 0 72.5 5 75.5 ;
      LAYER METS2 ;
        RECT 0 72.5 5 75.5 ;
      LAYER METS3 ;
        RECT 0 72.5 5 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 5 111.5 ;
      LAYER MET6 ;
        RECT 0 108.5 5 111.5 ;
      LAYER METG1 ;
        RECT 0 108.5 5 111.5 ;
      LAYER METS1 ;
        RECT 0 108.5 5 111.5 ;
      LAYER METS2 ;
        RECT 0 108.5 5 111.5 ;
      LAYER METS3 ;
        RECT 0 108.5 5 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 5 131.5 ;
      LAYER MET6 ;
        RECT 0 128.5 5 131.5 ;
      LAYER METG1 ;
        RECT 0 128.5 5 131.5 ;
      LAYER METS1 ;
        RECT 0 128.5 5 131.5 ;
      LAYER METS2 ;
        RECT 0 128.5 5 131.5 ;
      LAYER METS3 ;
        RECT 0 128.5 5 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 5 139.5 ;
      LAYER MET6 ;
        RECT 0 136.5 5 139.5 ;
      LAYER METG1 ;
        RECT 0 136.5 5 139.5 ;
      LAYER METS1 ;
        RECT 0 136.5 5 139.5 ;
      LAYER METS2 ;
        RECT 0 136.5 5 139.5 ;
      LAYER METS3 ;
        RECT 0 136.5 5 139.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 75.6 5 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 5 79.5 ;
      LAYER MET6 ;
        RECT 0 76.5 5 79.5 ;
      LAYER METG1 ;
        RECT 0 76.5 5 79.5 ;
      LAYER METS1 ;
        RECT 0 76.5 5 79.5 ;
      LAYER METS2 ;
        RECT 0 76.5 5 79.5 ;
      LAYER METS3 ;
        RECT 0 76.5 5 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 5 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 5 83.5 ;
      LAYER MET6 ;
        RECT 0 80.5 5 83.5 ;
      LAYER METG1 ;
        RECT 0 80.5 5 83.5 ;
      LAYER METS1 ;
        RECT 0 80.5 5 83.5 ;
      LAYER METS2 ;
        RECT 0 80.5 5 83.5 ;
      LAYER METS3 ;
        RECT 0 80.5 5 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 5 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 5 87.5 ;
      LAYER MET6 ;
        RECT 0 84.5 5 87.5 ;
      LAYER METG1 ;
        RECT 0 84.5 5 87.5 ;
      LAYER METS1 ;
        RECT 0 84.5 5 87.5 ;
      LAYER METS2 ;
        RECT 0 84.5 5 87.5 ;
      LAYER METS3 ;
        RECT 0 84.5 5 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 5 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 5 91.5 ;
      LAYER MET6 ;
        RECT 0 88.5 5 91.5 ;
      LAYER METG1 ;
        RECT 0 88.5 5 91.5 ;
      LAYER METS1 ;
        RECT 0 88.5 5 91.5 ;
      LAYER METS2 ;
        RECT 0 88.5 5 91.5 ;
      LAYER METS3 ;
        RECT 0 88.5 5 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 5 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 5 95.5 ;
      LAYER MET6 ;
        RECT 0 92.5 5 95.5 ;
      LAYER METG1 ;
        RECT 0 92.5 5 95.5 ;
      LAYER METS1 ;
        RECT 0 92.5 5 95.5 ;
      LAYER METS2 ;
        RECT 0 92.5 5 95.5 ;
      LAYER METS3 ;
        RECT 0 92.5 5 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 5 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 5 99.5 ;
      LAYER MET6 ;
        RECT 0 96.5 5 99.5 ;
      LAYER METG1 ;
        RECT 0 96.5 5 99.5 ;
      LAYER METS1 ;
        RECT 0 96.5 5 99.5 ;
      LAYER METS2 ;
        RECT 0 96.5 5 99.5 ;
      LAYER METS3 ;
        RECT 0 96.5 5 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 5 155.5 ;
      LAYER MET6 ;
        RECT 0 152.5 5 155.5 ;
      LAYER METG1 ;
        RECT 0 152.5 5 155.5 ;
      LAYER METS1 ;
        RECT 0 152.5 5 155.5 ;
      LAYER METS2 ;
        RECT 0 152.5 5 155.5 ;
      LAYER METS3 ;
        RECT 0 152.5 5 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 5 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 5 159.5 ;
      LAYER MET6 ;
        RECT 0 156.5 5 159.5 ;
      LAYER METG1 ;
        RECT 0 156.5 5 159.5 ;
      LAYER METS1 ;
        RECT 0 156.5 5 159.5 ;
      LAYER METS2 ;
        RECT 0 156.5 5 159.5 ;
      LAYER METS3 ;
        RECT 0 156.5 5 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 5 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 5 163.5 ;
      LAYER MET6 ;
        RECT 0 160.5 5 163.5 ;
      LAYER METG1 ;
        RECT 0 160.5 5 163.5 ;
      LAYER METS1 ;
        RECT 0 160.5 5 163.5 ;
      LAYER METS2 ;
        RECT 0 160.5 5 163.5 ;
      LAYER METS3 ;
        RECT 0 160.5 5 163.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 4.5 5 7.5 ;
      LAYER MET6 ;
        RECT 0 4.5 5 7.5 ;
      LAYER METG1 ;
        RECT 0 4.5 5 7.5 ;
      LAYER METS1 ;
        RECT 0 4.5 5 7.5 ;
      LAYER METS2 ;
        RECT 0 4.5 5 7.5 ;
      LAYER METS3 ;
        RECT 0 4.5 5 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 5 11.5 ;
      LAYER MET6 ;
        RECT 0 8.5 5 11.5 ;
      LAYER METG1 ;
        RECT 0 8.5 5 11.5 ;
      LAYER METS1 ;
        RECT 0 8.5 5 11.5 ;
      LAYER METS2 ;
        RECT 0 8.5 5 11.5 ;
      LAYER METS3 ;
        RECT 0 8.5 5 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 5 23.5 ;
      LAYER MET6 ;
        RECT 0 20.5 5 23.5 ;
      LAYER METG1 ;
        RECT 0 20.5 5 23.5 ;
      LAYER METS1 ;
        RECT 0 20.5 5 23.5 ;
      LAYER METS2 ;
        RECT 0 20.5 5 23.5 ;
      LAYER METS3 ;
        RECT 0 20.5 5 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 5 27.5 ;
      LAYER MET6 ;
        RECT 0 24.5 5 27.5 ;
      LAYER METG1 ;
        RECT 0 24.5 5 27.5 ;
      LAYER METS1 ;
        RECT 0 24.5 5 27.5 ;
      LAYER METS2 ;
        RECT 0 24.5 5 27.5 ;
      LAYER METS3 ;
        RECT 0 24.5 5 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 5 39.5 ;
      LAYER MET6 ;
        RECT 0 36.5 5 39.5 ;
      LAYER METG1 ;
        RECT 0 36.5 5 39.5 ;
      LAYER METS1 ;
        RECT 0 36.5 5 39.5 ;
      LAYER METS2 ;
        RECT 0 36.5 5 39.5 ;
      LAYER METS3 ;
        RECT 0 36.5 5 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 5 47.5 ;
      LAYER MET6 ;
        RECT 0 44.5 5 47.5 ;
      LAYER METG1 ;
        RECT 0 44.5 5 47.5 ;
      LAYER METS1 ;
        RECT 0 44.5 5 47.5 ;
      LAYER METS2 ;
        RECT 0 44.5 5 47.5 ;
      LAYER METS3 ;
        RECT 0 44.5 5 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 5 55.5 ;
      LAYER MET6 ;
        RECT 0 52.5 5 55.5 ;
      LAYER METG1 ;
        RECT 0 52.5 5 55.5 ;
      LAYER METS1 ;
        RECT 0 52.5 5 55.5 ;
      LAYER METS2 ;
        RECT 0 52.5 5 55.5 ;
      LAYER METS3 ;
        RECT 0 52.5 5 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 5 63.5 ;
      LAYER MET6 ;
        RECT 0 60.5 5 63.5 ;
      LAYER METG1 ;
        RECT 0 60.5 5 63.5 ;
      LAYER METS1 ;
        RECT 0 60.5 5 63.5 ;
      LAYER METS2 ;
        RECT 0 60.5 5 63.5 ;
      LAYER METS3 ;
        RECT 0 60.5 5 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 5 71.5 ;
      LAYER MET6 ;
        RECT 0 68.5 5 71.5 ;
      LAYER METG1 ;
        RECT 0 68.5 5 71.5 ;
      LAYER METS1 ;
        RECT 0 68.5 5 71.5 ;
      LAYER METS2 ;
        RECT 0 68.5 5 71.5 ;
      LAYER METS3 ;
        RECT 0 68.5 5 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 5 103.5 ;
      LAYER MET6 ;
        RECT 0 100.5 5 103.5 ;
      LAYER METG1 ;
        RECT 0 100.5 5 103.5 ;
      LAYER METS1 ;
        RECT 0 100.5 5 103.5 ;
      LAYER METS2 ;
        RECT 0 100.5 5 103.5 ;
      LAYER METS3 ;
        RECT 0 100.5 5 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 5 135.5 ;
      LAYER MET6 ;
        RECT 0 132.5 5 135.5 ;
      LAYER METG1 ;
        RECT 0 132.5 5 135.5 ;
      LAYER METS1 ;
        RECT 0 132.5 5 135.5 ;
      LAYER METS2 ;
        RECT 0 132.5 5 135.5 ;
      LAYER METS3 ;
        RECT 0 132.5 5 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 103.6 5 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 5 107.5 ;
      LAYER MET6 ;
        RECT 0 104.5 5 107.5 ;
      LAYER METG1 ;
        RECT 0 104.5 5 107.5 ;
      LAYER METS1 ;
        RECT 0 104.5 5 107.5 ;
      LAYER METS2 ;
        RECT 0 104.5 5 107.5 ;
      LAYER METS3 ;
        RECT 0 104.5 5 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 5 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 5 115.5 ;
      LAYER MET6 ;
        RECT 0 112.5 5 115.5 ;
      LAYER METG1 ;
        RECT 0 112.5 5 115.5 ;
      LAYER METS1 ;
        RECT 0 112.5 5 115.5 ;
      LAYER METS2 ;
        RECT 0 112.5 5 115.5 ;
      LAYER METS3 ;
        RECT 0 112.5 5 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 5 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 5 119.5 ;
      LAYER MET6 ;
        RECT 0 116.5 5 119.5 ;
      LAYER METG1 ;
        RECT 0 116.5 5 119.5 ;
      LAYER METS1 ;
        RECT 0 116.5 5 119.5 ;
      LAYER METS2 ;
        RECT 0 116.5 5 119.5 ;
      LAYER METS3 ;
        RECT 0 116.5 5 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 5 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 5 123.5 ;
      LAYER MET6 ;
        RECT 0 120.5 5 123.5 ;
      LAYER METG1 ;
        RECT 0 120.5 5 123.5 ;
      LAYER METS1 ;
        RECT 0 120.5 5 123.5 ;
      LAYER METS2 ;
        RECT 0 120.5 5 123.5 ;
      LAYER METS3 ;
        RECT 0 120.5 5 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 5 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 5 127.5 ;
      LAYER MET6 ;
        RECT 0 124.5 5 127.5 ;
      LAYER METG1 ;
        RECT 0 124.5 5 127.5 ;
      LAYER METS1 ;
        RECT 0 124.5 5 127.5 ;
      LAYER METS2 ;
        RECT 0 124.5 5 127.5 ;
      LAYER METS3 ;
        RECT 0 124.5 5 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 5 143.5 ;
      LAYER MET6 ;
        RECT 0 140.5 5 143.5 ;
      LAYER METG1 ;
        RECT 0 140.5 5 143.5 ;
      LAYER METS1 ;
        RECT 0 140.5 5 143.5 ;
      LAYER METS2 ;
        RECT 0 140.5 5 143.5 ;
      LAYER METS3 ;
        RECT 0 140.5 5 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 5 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 5 147.5 ;
      LAYER MET6 ;
        RECT 0 144.5 5 147.5 ;
      LAYER METG1 ;
        RECT 0 144.5 5 147.5 ;
      LAYER METS1 ;
        RECT 0 144.5 5 147.5 ;
      LAYER METS2 ;
        RECT 0 144.5 5 147.5 ;
      LAYER METS3 ;
        RECT 0 144.5 5 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 5 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 5 151.5 ;
      LAYER MET6 ;
        RECT 0 148.5 5 151.5 ;
      LAYER METG1 ;
        RECT 0 148.5 5 151.5 ;
      LAYER METS1 ;
        RECT 0 148.5 5 151.5 ;
      LAYER METS2 ;
        RECT 0 148.5 5 151.5 ;
      LAYER METS3 ;
        RECT 0 148.5 5 151.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 5 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 5 15.5 ;
      LAYER MET6 ;
        RECT 0 12.5 5 15.5 ;
      LAYER METG1 ;
        RECT 0 12.5 5 15.5 ;
      LAYER METS1 ;
        RECT 0 12.5 5 15.5 ;
      LAYER METS2 ;
        RECT 0 12.5 5 15.5 ;
      LAYER METS3 ;
        RECT 0 12.5 5 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 5 19.5 ;
      LAYER MET6 ;
        RECT 0 16.5 5 19.5 ;
      LAYER METG1 ;
        RECT 0 16.5 5 19.5 ;
      LAYER METS1 ;
        RECT 0 16.5 5 19.5 ;
      LAYER METS2 ;
        RECT 0 16.5 5 19.5 ;
      LAYER METS3 ;
        RECT 0 16.5 5 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 5 170 ;
    LAYER CUT12 ;
      RECT 0 0 5 170 ;
    LAYER MET2 ;
      RECT 0 0 5 170 ;
    LAYER CUT23 ;
      RECT 0 0 5 170 ;
    LAYER MET3 ;
      RECT 0 0 5 170 ;
    LAYER CUT34 ;
      RECT 0 0 5 170 ;
    LAYER MET4 ;
      RECT 0 0 5 170 ;
    LAYER CUT45 ;
      RECT 0 0 5 170 ;
    LAYER MET5 ;
      RECT 0 0 5 170 ;
    LAYER CUT56 ;
      RECT 0 0 5 170 ;
    LAYER MET6 ;
      RECT 0 0 5 170 ;
    LAYER CUTS1 ;
      RECT 0 0 5 170 ;
    LAYER METS1 ;
      RECT 0 0 5 170 ;
    LAYER CUTS2 ;
      RECT 0 0 5 170 ;
    LAYER METS2 ;
      RECT 0 0 5 170 ;
    LAYER CUTS3 ;
      RECT 0 0 5 170 ;
    LAYER METS3 ;
      RECT 0 0 5 170 ;
    LAYER CUTG1 ;
      RECT 0 0 5 170 ;
    LAYER METG1 ;
      RECT 0 0 5 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 5.000 2.000 ;
  END
END IOCB2ES54C0A1


MACRO IOCB2ESA4C0A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2ESA4C0A1 0 0 ;
  SIZE 10 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 28.5 10 31.5 ;
      LAYER MET6 ;
        RECT 0 28.5 10 31.5 ;
      LAYER METG1 ;
        RECT 0 28.5 10 31.5 ;
      LAYER METS1 ;
        RECT 0 28.5 10 31.5 ;
      LAYER METS2 ;
        RECT 0 28.5 10 31.5 ;
      LAYER METS3 ;
        RECT 0 28.5 10 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 10 35.5 ;
      LAYER MET6 ;
        RECT 0 32.5 10 35.5 ;
      LAYER METG1 ;
        RECT 0 32.5 10 35.5 ;
      LAYER METS1 ;
        RECT 0 32.5 10 35.5 ;
      LAYER METS2 ;
        RECT 0 32.5 10 35.5 ;
      LAYER METS3 ;
        RECT 0 32.5 10 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 10 43.5 ;
      LAYER MET6 ;
        RECT 0 40.5 10 43.5 ;
      LAYER METG1 ;
        RECT 0 40.5 10 43.5 ;
      LAYER METS1 ;
        RECT 0 40.5 10 43.5 ;
      LAYER METS2 ;
        RECT 0 40.5 10 43.5 ;
      LAYER METS3 ;
        RECT 0 40.5 10 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 10 51.5 ;
      LAYER MET6 ;
        RECT 0 48.5 10 51.5 ;
      LAYER METG1 ;
        RECT 0 48.5 10 51.5 ;
      LAYER METS1 ;
        RECT 0 48.5 10 51.5 ;
      LAYER METS2 ;
        RECT 0 48.5 10 51.5 ;
      LAYER METS3 ;
        RECT 0 48.5 10 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 10 59.5 ;
      LAYER MET6 ;
        RECT 0 56.5 10 59.5 ;
      LAYER METG1 ;
        RECT 0 56.5 10 59.5 ;
      LAYER METS1 ;
        RECT 0 56.5 10 59.5 ;
      LAYER METS2 ;
        RECT 0 56.5 10 59.5 ;
      LAYER METS3 ;
        RECT 0 56.5 10 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 10 67.5 ;
      LAYER MET6 ;
        RECT 0 64.5 10 67.5 ;
      LAYER METG1 ;
        RECT 0 64.5 10 67.5 ;
      LAYER METS1 ;
        RECT 0 64.5 10 67.5 ;
      LAYER METS2 ;
        RECT 0 64.5 10 67.5 ;
      LAYER METS3 ;
        RECT 0 64.5 10 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 10 75.5 ;
      LAYER MET6 ;
        RECT 0 72.5 10 75.5 ;
      LAYER METG1 ;
        RECT 0 72.5 10 75.5 ;
      LAYER METS1 ;
        RECT 0 72.5 10 75.5 ;
      LAYER METS2 ;
        RECT 0 72.5 10 75.5 ;
      LAYER METS3 ;
        RECT 0 72.5 10 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 10 111.5 ;
      LAYER MET6 ;
        RECT 0 108.5 10 111.5 ;
      LAYER METG1 ;
        RECT 0 108.5 10 111.5 ;
      LAYER METS1 ;
        RECT 0 108.5 10 111.5 ;
      LAYER METS2 ;
        RECT 0 108.5 10 111.5 ;
      LAYER METS3 ;
        RECT 0 108.5 10 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 10 131.5 ;
      LAYER MET6 ;
        RECT 0 128.5 10 131.5 ;
      LAYER METG1 ;
        RECT 0 128.5 10 131.5 ;
      LAYER METS1 ;
        RECT 0 128.5 10 131.5 ;
      LAYER METS2 ;
        RECT 0 128.5 10 131.5 ;
      LAYER METS3 ;
        RECT 0 128.5 10 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 10 139.5 ;
      LAYER MET6 ;
        RECT 0 136.5 10 139.5 ;
      LAYER METG1 ;
        RECT 0 136.5 10 139.5 ;
      LAYER METS1 ;
        RECT 0 136.5 10 139.5 ;
      LAYER METS2 ;
        RECT 0 136.5 10 139.5 ;
      LAYER METS3 ;
        RECT 0 136.5 10 139.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 75.6 10 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 10 79.5 ;
      LAYER MET6 ;
        RECT 0 76.5 10 79.5 ;
      LAYER METG1 ;
        RECT 0 76.5 10 79.5 ;
      LAYER METS1 ;
        RECT 0 76.5 10 79.5 ;
      LAYER METS2 ;
        RECT 0 76.5 10 79.5 ;
      LAYER METS3 ;
        RECT 0 76.5 10 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 10 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 10 83.5 ;
      LAYER MET6 ;
        RECT 0 80.5 10 83.5 ;
      LAYER METG1 ;
        RECT 0 80.5 10 83.5 ;
      LAYER METS1 ;
        RECT 0 80.5 10 83.5 ;
      LAYER METS2 ;
        RECT 0 80.5 10 83.5 ;
      LAYER METS3 ;
        RECT 0 80.5 10 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 10 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 10 87.5 ;
      LAYER MET6 ;
        RECT 0 84.5 10 87.5 ;
      LAYER METG1 ;
        RECT 0 84.5 10 87.5 ;
      LAYER METS1 ;
        RECT 0 84.5 10 87.5 ;
      LAYER METS2 ;
        RECT 0 84.5 10 87.5 ;
      LAYER METS3 ;
        RECT 0 84.5 10 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 10 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 10 91.5 ;
      LAYER MET6 ;
        RECT 0 88.5 10 91.5 ;
      LAYER METG1 ;
        RECT 0 88.5 10 91.5 ;
      LAYER METS1 ;
        RECT 0 88.5 10 91.5 ;
      LAYER METS2 ;
        RECT 0 88.5 10 91.5 ;
      LAYER METS3 ;
        RECT 0 88.5 10 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 10 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 10 95.5 ;
      LAYER MET6 ;
        RECT 0 92.5 10 95.5 ;
      LAYER METG1 ;
        RECT 0 92.5 10 95.5 ;
      LAYER METS1 ;
        RECT 0 92.5 10 95.5 ;
      LAYER METS2 ;
        RECT 0 92.5 10 95.5 ;
      LAYER METS3 ;
        RECT 0 92.5 10 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 10 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 10 99.5 ;
      LAYER MET6 ;
        RECT 0 96.5 10 99.5 ;
      LAYER METG1 ;
        RECT 0 96.5 10 99.5 ;
      LAYER METS1 ;
        RECT 0 96.5 10 99.5 ;
      LAYER METS2 ;
        RECT 0 96.5 10 99.5 ;
      LAYER METS3 ;
        RECT 0 96.5 10 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 10 155.5 ;
      LAYER MET6 ;
        RECT 0 152.5 10 155.5 ;
      LAYER METG1 ;
        RECT 0 152.5 10 155.5 ;
      LAYER METS1 ;
        RECT 0 152.5 10 155.5 ;
      LAYER METS2 ;
        RECT 0 152.5 10 155.5 ;
      LAYER METS3 ;
        RECT 0 152.5 10 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 10 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 10 159.5 ;
      LAYER MET6 ;
        RECT 0 156.5 10 159.5 ;
      LAYER METG1 ;
        RECT 0 156.5 10 159.5 ;
      LAYER METS1 ;
        RECT 0 156.5 10 159.5 ;
      LAYER METS2 ;
        RECT 0 156.5 10 159.5 ;
      LAYER METS3 ;
        RECT 0 156.5 10 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 10 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 10 163.5 ;
      LAYER MET6 ;
        RECT 0 160.5 10 163.5 ;
      LAYER METG1 ;
        RECT 0 160.5 10 163.5 ;
      LAYER METS1 ;
        RECT 0 160.5 10 163.5 ;
      LAYER METS2 ;
        RECT 0 160.5 10 163.5 ;
      LAYER METS3 ;
        RECT 0 160.5 10 163.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 4.5 10 7.5 ;
      LAYER MET6 ;
        RECT 0 4.5 10 7.5 ;
      LAYER METG1 ;
        RECT 0 4.5 10 7.5 ;
      LAYER METS1 ;
        RECT 0 4.5 10 7.5 ;
      LAYER METS2 ;
        RECT 0 4.5 10 7.5 ;
      LAYER METS3 ;
        RECT 0 4.5 10 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 10 11.5 ;
      LAYER MET6 ;
        RECT 0 8.5 10 11.5 ;
      LAYER METG1 ;
        RECT 0 8.5 10 11.5 ;
      LAYER METS1 ;
        RECT 0 8.5 10 11.5 ;
      LAYER METS2 ;
        RECT 0 8.5 10 11.5 ;
      LAYER METS3 ;
        RECT 0 8.5 10 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 10 23.5 ;
      LAYER MET6 ;
        RECT 0 20.5 10 23.5 ;
      LAYER METG1 ;
        RECT 0 20.5 10 23.5 ;
      LAYER METS1 ;
        RECT 0 20.5 10 23.5 ;
      LAYER METS2 ;
        RECT 0 20.5 10 23.5 ;
      LAYER METS3 ;
        RECT 0 20.5 10 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 10 27.5 ;
      LAYER MET6 ;
        RECT 0 24.5 10 27.5 ;
      LAYER METG1 ;
        RECT 0 24.5 10 27.5 ;
      LAYER METS1 ;
        RECT 0 24.5 10 27.5 ;
      LAYER METS2 ;
        RECT 0 24.5 10 27.5 ;
      LAYER METS3 ;
        RECT 0 24.5 10 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 10 39.5 ;
      LAYER MET6 ;
        RECT 0 36.5 10 39.5 ;
      LAYER METG1 ;
        RECT 0 36.5 10 39.5 ;
      LAYER METS1 ;
        RECT 0 36.5 10 39.5 ;
      LAYER METS2 ;
        RECT 0 36.5 10 39.5 ;
      LAYER METS3 ;
        RECT 0 36.5 10 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 10 47.5 ;
      LAYER MET6 ;
        RECT 0 44.5 10 47.5 ;
      LAYER METG1 ;
        RECT 0 44.5 10 47.5 ;
      LAYER METS1 ;
        RECT 0 44.5 10 47.5 ;
      LAYER METS2 ;
        RECT 0 44.5 10 47.5 ;
      LAYER METS3 ;
        RECT 0 44.5 10 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 10 55.5 ;
      LAYER MET6 ;
        RECT 0 52.5 10 55.5 ;
      LAYER METG1 ;
        RECT 0 52.5 10 55.5 ;
      LAYER METS1 ;
        RECT 0 52.5 10 55.5 ;
      LAYER METS2 ;
        RECT 0 52.5 10 55.5 ;
      LAYER METS3 ;
        RECT 0 52.5 10 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 10 63.5 ;
      LAYER MET6 ;
        RECT 0 60.5 10 63.5 ;
      LAYER METG1 ;
        RECT 0 60.5 10 63.5 ;
      LAYER METS1 ;
        RECT 0 60.5 10 63.5 ;
      LAYER METS2 ;
        RECT 0 60.5 10 63.5 ;
      LAYER METS3 ;
        RECT 0 60.5 10 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 10 71.5 ;
      LAYER MET6 ;
        RECT 0 68.5 10 71.5 ;
      LAYER METG1 ;
        RECT 0 68.5 10 71.5 ;
      LAYER METS1 ;
        RECT 0 68.5 10 71.5 ;
      LAYER METS2 ;
        RECT 0 68.5 10 71.5 ;
      LAYER METS3 ;
        RECT 0 68.5 10 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 10 103.5 ;
      LAYER MET6 ;
        RECT 0 100.5 10 103.5 ;
      LAYER METG1 ;
        RECT 0 100.5 10 103.5 ;
      LAYER METS1 ;
        RECT 0 100.5 10 103.5 ;
      LAYER METS2 ;
        RECT 0 100.5 10 103.5 ;
      LAYER METS3 ;
        RECT 0 100.5 10 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 10 135.5 ;
      LAYER MET6 ;
        RECT 0 132.5 10 135.5 ;
      LAYER METG1 ;
        RECT 0 132.5 10 135.5 ;
      LAYER METS1 ;
        RECT 0 132.5 10 135.5 ;
      LAYER METS2 ;
        RECT 0 132.5 10 135.5 ;
      LAYER METS3 ;
        RECT 0 132.5 10 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 103.6 10 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 10 107.5 ;
      LAYER MET6 ;
        RECT 0 104.5 10 107.5 ;
      LAYER METG1 ;
        RECT 0 104.5 10 107.5 ;
      LAYER METS1 ;
        RECT 0 104.5 10 107.5 ;
      LAYER METS2 ;
        RECT 0 104.5 10 107.5 ;
      LAYER METS3 ;
        RECT 0 104.5 10 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 10 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 10 115.5 ;
      LAYER MET6 ;
        RECT 0 112.5 10 115.5 ;
      LAYER METG1 ;
        RECT 0 112.5 10 115.5 ;
      LAYER METS1 ;
        RECT 0 112.5 10 115.5 ;
      LAYER METS2 ;
        RECT 0 112.5 10 115.5 ;
      LAYER METS3 ;
        RECT 0 112.5 10 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 10 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 10 119.5 ;
      LAYER MET6 ;
        RECT 0 116.5 10 119.5 ;
      LAYER METG1 ;
        RECT 0 116.5 10 119.5 ;
      LAYER METS1 ;
        RECT 0 116.5 10 119.5 ;
      LAYER METS2 ;
        RECT 0 116.5 10 119.5 ;
      LAYER METS3 ;
        RECT 0 116.5 10 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 10 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 10 123.5 ;
      LAYER MET6 ;
        RECT 0 120.5 10 123.5 ;
      LAYER METG1 ;
        RECT 0 120.5 10 123.5 ;
      LAYER METS1 ;
        RECT 0 120.5 10 123.5 ;
      LAYER METS2 ;
        RECT 0 120.5 10 123.5 ;
      LAYER METS3 ;
        RECT 0 120.5 10 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 10 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 10 127.5 ;
      LAYER MET6 ;
        RECT 0 124.5 10 127.5 ;
      LAYER METG1 ;
        RECT 0 124.5 10 127.5 ;
      LAYER METS1 ;
        RECT 0 124.5 10 127.5 ;
      LAYER METS2 ;
        RECT 0 124.5 10 127.5 ;
      LAYER METS3 ;
        RECT 0 124.5 10 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 10 143.5 ;
      LAYER MET6 ;
        RECT 0 140.5 10 143.5 ;
      LAYER METG1 ;
        RECT 0 140.5 10 143.5 ;
      LAYER METS1 ;
        RECT 0 140.5 10 143.5 ;
      LAYER METS2 ;
        RECT 0 140.5 10 143.5 ;
      LAYER METS3 ;
        RECT 0 140.5 10 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 10 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 10 147.5 ;
      LAYER MET6 ;
        RECT 0 144.5 10 147.5 ;
      LAYER METG1 ;
        RECT 0 144.5 10 147.5 ;
      LAYER METS1 ;
        RECT 0 144.5 10 147.5 ;
      LAYER METS2 ;
        RECT 0 144.5 10 147.5 ;
      LAYER METS3 ;
        RECT 0 144.5 10 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 10 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 10 151.5 ;
      LAYER MET6 ;
        RECT 0 148.5 10 151.5 ;
      LAYER METG1 ;
        RECT 0 148.5 10 151.5 ;
      LAYER METS1 ;
        RECT 0 148.5 10 151.5 ;
      LAYER METS2 ;
        RECT 0 148.5 10 151.5 ;
      LAYER METS3 ;
        RECT 0 148.5 10 151.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 10 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 10 15.5 ;
      LAYER MET6 ;
        RECT 0 12.5 10 15.5 ;
      LAYER METG1 ;
        RECT 0 12.5 10 15.5 ;
      LAYER METS1 ;
        RECT 0 12.5 10 15.5 ;
      LAYER METS2 ;
        RECT 0 12.5 10 15.5 ;
      LAYER METS3 ;
        RECT 0 12.5 10 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 10 19.5 ;
      LAYER MET6 ;
        RECT 0 16.5 10 19.5 ;
      LAYER METG1 ;
        RECT 0 16.5 10 19.5 ;
      LAYER METS1 ;
        RECT 0 16.5 10 19.5 ;
      LAYER METS2 ;
        RECT 0 16.5 10 19.5 ;
      LAYER METS3 ;
        RECT 0 16.5 10 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 10 170 ;
    LAYER CUT12 ;
      RECT 0 0 10 170 ;
    LAYER MET2 ;
      RECT 0 0 10 170 ;
    LAYER CUT23 ;
      RECT 0 0 10 170 ;
    LAYER MET3 ;
      RECT 0 0 10 170 ;
    LAYER CUT34 ;
      RECT 0 0 10 170 ;
    LAYER MET4 ;
      RECT 0 0 10 170 ;
    LAYER CUT45 ;
      RECT 0 0 10 170 ;
    LAYER MET5 ;
      RECT 0 0 10 170 ;
    LAYER CUT56 ;
      RECT 0 0 10 170 ;
    LAYER MET6 ;
      RECT 0 0 10 170 ;
    LAYER CUTS1 ;
      RECT 0 0 10 170 ;
    LAYER METS1 ;
      RECT 0 0 10 170 ;
    LAYER CUTS2 ;
      RECT 0 0 10 170 ;
    LAYER METS2 ;
      RECT 0 0 10 170 ;
    LAYER CUTS3 ;
      RECT 0 0 10 170 ;
    LAYER METS3 ;
      RECT 0 0 10 170 ;
    LAYER CUTG1 ;
      RECT 0 0 10 170 ;
    LAYER METG1 ;
      RECT 0 0 10 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 10.000 2.000 ;
  END
END IOCB2ESA4C0A1


MACRO IOCB2ESB4C0A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2ESB4C0A1 0 0 ;
  SIZE 0.1 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 28.5 0.1 31.5 ;
      LAYER MET6 ;
        RECT 0 28.5 0.1 31.5 ;
      LAYER METG1 ;
        RECT 0 28.5 0.1 31.5 ;
      LAYER METS1 ;
        RECT 0 28.5 0.1 31.5 ;
      LAYER METS2 ;
        RECT 0 28.5 0.1 31.5 ;
      LAYER METS3 ;
        RECT 0 28.5 0.1 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 0.1 35.5 ;
      LAYER MET6 ;
        RECT 0 32.5 0.1 35.5 ;
      LAYER METG1 ;
        RECT 0 32.5 0.1 35.5 ;
      LAYER METS1 ;
        RECT 0 32.5 0.1 35.5 ;
      LAYER METS2 ;
        RECT 0 32.5 0.1 35.5 ;
      LAYER METS3 ;
        RECT 0 32.5 0.1 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 0.1 43.5 ;
      LAYER MET6 ;
        RECT 0 40.5 0.1 43.5 ;
      LAYER METG1 ;
        RECT 0 40.5 0.1 43.5 ;
      LAYER METS1 ;
        RECT 0 40.5 0.1 43.5 ;
      LAYER METS2 ;
        RECT 0 40.5 0.1 43.5 ;
      LAYER METS3 ;
        RECT 0 40.5 0.1 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 0.1 51.5 ;
      LAYER MET6 ;
        RECT 0 48.5 0.1 51.5 ;
      LAYER METG1 ;
        RECT 0 48.5 0.1 51.5 ;
      LAYER METS1 ;
        RECT 0 48.5 0.1 51.5 ;
      LAYER METS2 ;
        RECT 0 48.5 0.1 51.5 ;
      LAYER METS3 ;
        RECT 0 48.5 0.1 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 0.1 59.5 ;
      LAYER MET6 ;
        RECT 0 56.5 0.1 59.5 ;
      LAYER METG1 ;
        RECT 0 56.5 0.1 59.5 ;
      LAYER METS1 ;
        RECT 0 56.5 0.1 59.5 ;
      LAYER METS2 ;
        RECT 0 56.5 0.1 59.5 ;
      LAYER METS3 ;
        RECT 0 56.5 0.1 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 0.1 67.5 ;
      LAYER MET6 ;
        RECT 0 64.5 0.1 67.5 ;
      LAYER METG1 ;
        RECT 0 64.5 0.1 67.5 ;
      LAYER METS1 ;
        RECT 0 64.5 0.1 67.5 ;
      LAYER METS2 ;
        RECT 0 64.5 0.1 67.5 ;
      LAYER METS3 ;
        RECT 0 64.5 0.1 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 0.1 75.5 ;
      LAYER MET6 ;
        RECT 0 72.5 0.1 75.5 ;
      LAYER METG1 ;
        RECT 0 72.5 0.1 75.5 ;
      LAYER METS1 ;
        RECT 0 72.5 0.1 75.5 ;
      LAYER METS2 ;
        RECT 0 72.5 0.1 75.5 ;
      LAYER METS3 ;
        RECT 0 72.5 0.1 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 0.1 111.5 ;
      LAYER MET6 ;
        RECT 0 108.5 0.1 111.5 ;
      LAYER METG1 ;
        RECT 0 108.5 0.1 111.5 ;
      LAYER METS1 ;
        RECT 0 108.5 0.1 111.5 ;
      LAYER METS2 ;
        RECT 0 108.5 0.1 111.5 ;
      LAYER METS3 ;
        RECT 0 108.5 0.1 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 0.1 131.5 ;
      LAYER MET6 ;
        RECT 0 128.5 0.1 131.5 ;
      LAYER METG1 ;
        RECT 0 128.5 0.1 131.5 ;
      LAYER METS1 ;
        RECT 0 128.5 0.1 131.5 ;
      LAYER METS2 ;
        RECT 0 128.5 0.1 131.5 ;
      LAYER METS3 ;
        RECT 0 128.5 0.1 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 0.1 139.5 ;
      LAYER MET6 ;
        RECT 0 136.5 0.1 139.5 ;
      LAYER METG1 ;
        RECT 0 136.5 0.1 139.5 ;
      LAYER METS1 ;
        RECT 0 136.5 0.1 139.5 ;
      LAYER METS2 ;
        RECT 0 136.5 0.1 139.5 ;
      LAYER METS3 ;
        RECT 0 136.5 0.1 139.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 75.6 0.1 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 0.1 79.5 ;
      LAYER MET6 ;
        RECT 0 76.5 0.1 79.5 ;
      LAYER METG1 ;
        RECT 0 76.5 0.1 79.5 ;
      LAYER METS1 ;
        RECT 0 76.5 0.1 79.5 ;
      LAYER METS2 ;
        RECT 0 76.5 0.1 79.5 ;
      LAYER METS3 ;
        RECT 0 76.5 0.1 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 0.1 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 0.1 83.5 ;
      LAYER MET6 ;
        RECT 0 80.5 0.1 83.5 ;
      LAYER METG1 ;
        RECT 0 80.5 0.1 83.5 ;
      LAYER METS1 ;
        RECT 0 80.5 0.1 83.5 ;
      LAYER METS2 ;
        RECT 0 80.5 0.1 83.5 ;
      LAYER METS3 ;
        RECT 0 80.5 0.1 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 0.1 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 0.1 87.5 ;
      LAYER MET6 ;
        RECT 0 84.5 0.1 87.5 ;
      LAYER METG1 ;
        RECT 0 84.5 0.1 87.5 ;
      LAYER METS1 ;
        RECT 0 84.5 0.1 87.5 ;
      LAYER METS2 ;
        RECT 0 84.5 0.1 87.5 ;
      LAYER METS3 ;
        RECT 0 84.5 0.1 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 0.1 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 0.1 91.5 ;
      LAYER MET6 ;
        RECT 0 88.5 0.1 91.5 ;
      LAYER METG1 ;
        RECT 0 88.5 0.1 91.5 ;
      LAYER METS1 ;
        RECT 0 88.5 0.1 91.5 ;
      LAYER METS2 ;
        RECT 0 88.5 0.1 91.5 ;
      LAYER METS3 ;
        RECT 0 88.5 0.1 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 0.1 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 0.1 95.5 ;
      LAYER MET6 ;
        RECT 0 92.5 0.1 95.5 ;
      LAYER METG1 ;
        RECT 0 92.5 0.1 95.5 ;
      LAYER METS1 ;
        RECT 0 92.5 0.1 95.5 ;
      LAYER METS2 ;
        RECT 0 92.5 0.1 95.5 ;
      LAYER METS3 ;
        RECT 0 92.5 0.1 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 0.1 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 0.1 99.5 ;
      LAYER MET6 ;
        RECT 0 96.5 0.1 99.5 ;
      LAYER METG1 ;
        RECT 0 96.5 0.1 99.5 ;
      LAYER METS1 ;
        RECT 0 96.5 0.1 99.5 ;
      LAYER METS2 ;
        RECT 0 96.5 0.1 99.5 ;
      LAYER METS3 ;
        RECT 0 96.5 0.1 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 0.1 155.5 ;
      LAYER MET6 ;
        RECT 0 152.5 0.1 155.5 ;
      LAYER METG1 ;
        RECT 0 152.5 0.1 155.5 ;
      LAYER METS1 ;
        RECT 0 152.5 0.1 155.5 ;
      LAYER METS2 ;
        RECT 0 152.5 0.1 155.5 ;
      LAYER METS3 ;
        RECT 0 152.5 0.1 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 0.1 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 0.1 159.5 ;
      LAYER MET6 ;
        RECT 0 156.5 0.1 159.5 ;
      LAYER METG1 ;
        RECT 0 156.5 0.1 159.5 ;
      LAYER METS1 ;
        RECT 0 156.5 0.1 159.5 ;
      LAYER METS2 ;
        RECT 0 156.5 0.1 159.5 ;
      LAYER METS3 ;
        RECT 0 156.5 0.1 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 0.1 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 0.1 163.5 ;
      LAYER MET6 ;
        RECT 0 160.5 0.1 163.5 ;
      LAYER METG1 ;
        RECT 0 160.5 0.1 163.5 ;
      LAYER METS1 ;
        RECT 0 160.5 0.1 163.5 ;
      LAYER METS2 ;
        RECT 0 160.5 0.1 163.5 ;
      LAYER METS3 ;
        RECT 0 160.5 0.1 163.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 4.5 0.1 7.5 ;
      LAYER MET6 ;
        RECT 0 4.5 0.1 7.5 ;
      LAYER METG1 ;
        RECT 0 4.5 0.1 7.5 ;
      LAYER METS1 ;
        RECT 0 4.5 0.1 7.5 ;
      LAYER METS2 ;
        RECT 0 4.5 0.1 7.5 ;
      LAYER METS3 ;
        RECT 0 4.5 0.1 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 0.1 11.5 ;
      LAYER MET6 ;
        RECT 0 8.5 0.1 11.5 ;
      LAYER METG1 ;
        RECT 0 8.5 0.1 11.5 ;
      LAYER METS1 ;
        RECT 0 8.5 0.1 11.5 ;
      LAYER METS2 ;
        RECT 0 8.5 0.1 11.5 ;
      LAYER METS3 ;
        RECT 0 8.5 0.1 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 0.1 23.5 ;
      LAYER MET6 ;
        RECT 0 20.5 0.1 23.5 ;
      LAYER METG1 ;
        RECT 0 20.5 0.1 23.5 ;
      LAYER METS1 ;
        RECT 0 20.5 0.1 23.5 ;
      LAYER METS2 ;
        RECT 0 20.5 0.1 23.5 ;
      LAYER METS3 ;
        RECT 0 20.5 0.1 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 0.1 27.5 ;
      LAYER MET6 ;
        RECT 0 24.5 0.1 27.5 ;
      LAYER METG1 ;
        RECT 0 24.5 0.1 27.5 ;
      LAYER METS1 ;
        RECT 0 24.5 0.1 27.5 ;
      LAYER METS2 ;
        RECT 0 24.5 0.1 27.5 ;
      LAYER METS3 ;
        RECT 0 24.5 0.1 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 0.1 39.5 ;
      LAYER MET6 ;
        RECT 0 36.5 0.1 39.5 ;
      LAYER METG1 ;
        RECT 0 36.5 0.1 39.5 ;
      LAYER METS1 ;
        RECT 0 36.5 0.1 39.5 ;
      LAYER METS2 ;
        RECT 0 36.5 0.1 39.5 ;
      LAYER METS3 ;
        RECT 0 36.5 0.1 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 0.1 47.5 ;
      LAYER MET6 ;
        RECT 0 44.5 0.1 47.5 ;
      LAYER METG1 ;
        RECT 0 44.5 0.1 47.5 ;
      LAYER METS1 ;
        RECT 0 44.5 0.1 47.5 ;
      LAYER METS2 ;
        RECT 0 44.5 0.1 47.5 ;
      LAYER METS3 ;
        RECT 0 44.5 0.1 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 0.1 55.5 ;
      LAYER MET6 ;
        RECT 0 52.5 0.1 55.5 ;
      LAYER METG1 ;
        RECT 0 52.5 0.1 55.5 ;
      LAYER METS1 ;
        RECT 0 52.5 0.1 55.5 ;
      LAYER METS2 ;
        RECT 0 52.5 0.1 55.5 ;
      LAYER METS3 ;
        RECT 0 52.5 0.1 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 0.1 63.5 ;
      LAYER MET6 ;
        RECT 0 60.5 0.1 63.5 ;
      LAYER METG1 ;
        RECT 0 60.5 0.1 63.5 ;
      LAYER METS1 ;
        RECT 0 60.5 0.1 63.5 ;
      LAYER METS2 ;
        RECT 0 60.5 0.1 63.5 ;
      LAYER METS3 ;
        RECT 0 60.5 0.1 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 0.1 71.5 ;
      LAYER MET6 ;
        RECT 0 68.5 0.1 71.5 ;
      LAYER METG1 ;
        RECT 0 68.5 0.1 71.5 ;
      LAYER METS1 ;
        RECT 0 68.5 0.1 71.5 ;
      LAYER METS2 ;
        RECT 0 68.5 0.1 71.5 ;
      LAYER METS3 ;
        RECT 0 68.5 0.1 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 0.1 103.5 ;
      LAYER MET6 ;
        RECT 0 100.5 0.1 103.5 ;
      LAYER METG1 ;
        RECT 0 100.5 0.1 103.5 ;
      LAYER METS1 ;
        RECT 0 100.5 0.1 103.5 ;
      LAYER METS2 ;
        RECT 0 100.5 0.1 103.5 ;
      LAYER METS3 ;
        RECT 0 100.5 0.1 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 0.1 135.5 ;
      LAYER MET6 ;
        RECT 0 132.5 0.1 135.5 ;
      LAYER METG1 ;
        RECT 0 132.5 0.1 135.5 ;
      LAYER METS1 ;
        RECT 0 132.5 0.1 135.5 ;
      LAYER METS2 ;
        RECT 0 132.5 0.1 135.5 ;
      LAYER METS3 ;
        RECT 0 132.5 0.1 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 103.6 0.1 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 0.1 107.5 ;
      LAYER MET6 ;
        RECT 0 104.5 0.1 107.5 ;
      LAYER METG1 ;
        RECT 0 104.5 0.1 107.5 ;
      LAYER METS1 ;
        RECT 0 104.5 0.1 107.5 ;
      LAYER METS2 ;
        RECT 0 104.5 0.1 107.5 ;
      LAYER METS3 ;
        RECT 0 104.5 0.1 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 0.1 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 0.1 115.5 ;
      LAYER MET6 ;
        RECT 0 112.5 0.1 115.5 ;
      LAYER METG1 ;
        RECT 0 112.5 0.1 115.5 ;
      LAYER METS1 ;
        RECT 0 112.5 0.1 115.5 ;
      LAYER METS2 ;
        RECT 0 112.5 0.1 115.5 ;
      LAYER METS3 ;
        RECT 0 112.5 0.1 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 0.1 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 0.1 119.5 ;
      LAYER MET6 ;
        RECT 0 116.5 0.1 119.5 ;
      LAYER METG1 ;
        RECT 0 116.5 0.1 119.5 ;
      LAYER METS1 ;
        RECT 0 116.5 0.1 119.5 ;
      LAYER METS2 ;
        RECT 0 116.5 0.1 119.5 ;
      LAYER METS3 ;
        RECT 0 116.5 0.1 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 0.1 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 0.1 123.5 ;
      LAYER MET6 ;
        RECT 0 120.5 0.1 123.5 ;
      LAYER METG1 ;
        RECT 0 120.5 0.1 123.5 ;
      LAYER METS1 ;
        RECT 0 120.5 0.1 123.5 ;
      LAYER METS2 ;
        RECT 0 120.5 0.1 123.5 ;
      LAYER METS3 ;
        RECT 0 120.5 0.1 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 0.1 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 0.1 127.5 ;
      LAYER MET6 ;
        RECT 0 124.5 0.1 127.5 ;
      LAYER METG1 ;
        RECT 0 124.5 0.1 127.5 ;
      LAYER METS1 ;
        RECT 0 124.5 0.1 127.5 ;
      LAYER METS2 ;
        RECT 0 124.5 0.1 127.5 ;
      LAYER METS3 ;
        RECT 0 124.5 0.1 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 0.1 143.5 ;
      LAYER MET6 ;
        RECT 0 140.5 0.1 143.5 ;
      LAYER METG1 ;
        RECT 0 140.5 0.1 143.5 ;
      LAYER METS1 ;
        RECT 0 140.5 0.1 143.5 ;
      LAYER METS2 ;
        RECT 0 140.5 0.1 143.5 ;
      LAYER METS3 ;
        RECT 0 140.5 0.1 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 0.1 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 0.1 147.5 ;
      LAYER MET6 ;
        RECT 0 144.5 0.1 147.5 ;
      LAYER METG1 ;
        RECT 0 144.5 0.1 147.5 ;
      LAYER METS1 ;
        RECT 0 144.5 0.1 147.5 ;
      LAYER METS2 ;
        RECT 0 144.5 0.1 147.5 ;
      LAYER METS3 ;
        RECT 0 144.5 0.1 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 0.1 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 0.1 151.5 ;
      LAYER MET6 ;
        RECT 0 148.5 0.1 151.5 ;
      LAYER METG1 ;
        RECT 0 148.5 0.1 151.5 ;
      LAYER METS1 ;
        RECT 0 148.5 0.1 151.5 ;
      LAYER METS2 ;
        RECT 0 148.5 0.1 151.5 ;
      LAYER METS3 ;
        RECT 0 148.5 0.1 151.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 0.1 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 0.1 15.5 ;
      LAYER MET6 ;
        RECT 0 12.5 0.1 15.5 ;
      LAYER METG1 ;
        RECT 0 12.5 0.1 15.5 ;
      LAYER METS1 ;
        RECT 0 12.5 0.1 15.5 ;
      LAYER METS2 ;
        RECT 0 12.5 0.1 15.5 ;
      LAYER METS3 ;
        RECT 0 12.5 0.1 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 0.1 19.5 ;
      LAYER MET6 ;
        RECT 0 16.5 0.1 19.5 ;
      LAYER METG1 ;
        RECT 0 16.5 0.1 19.5 ;
      LAYER METS1 ;
        RECT 0 16.5 0.1 19.5 ;
      LAYER METS2 ;
        RECT 0 16.5 0.1 19.5 ;
      LAYER METS3 ;
        RECT 0 16.5 0.1 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 0.1 170 ;
    LAYER CUT12 ;
      RECT 0 0 0.1 170 ;
    LAYER MET2 ;
      RECT 0 0 0.1 170 ;
    LAYER CUT23 ;
      RECT 0 0 0.1 170 ;
    LAYER MET3 ;
      RECT 0 0 0.1 170 ;
    LAYER CUT34 ;
      RECT 0 0 0.1 170 ;
    LAYER MET4 ;
      RECT 0 0 0.1 170 ;
    LAYER CUT45 ;
      RECT 0 0 0.1 170 ;
    LAYER MET5 ;
      RECT 0 0 0.1 170 ;
    LAYER CUT56 ;
      RECT 0 0 0.1 170 ;
    LAYER MET6 ;
      RECT 0 0 0.1 170 ;
    LAYER CUTS1 ;
      RECT 0 0 0.1 170 ;
    LAYER METS1 ;
      RECT 0 0 0.1 170 ;
    LAYER CUTS2 ;
      RECT 0 0 0.1 170 ;
    LAYER METS2 ;
      RECT 0 0 0.1 170 ;
    LAYER CUTS3 ;
      RECT 0 0 0.1 170 ;
    LAYER METS3 ;
      RECT 0 0 0.1 170 ;
    LAYER CUTG1 ;
      RECT 0 0 0.1 170 ;
    LAYER METG1 ;
      RECT 0 0 0.1 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 0.100 2.000 ;
  END
END IOCB2ESB4C0A1


MACRO IOCB2ESD4C0A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2ESD4C0A1 0 0 ;
  SIZE 20 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 28.5 20 31.5 ;
      LAYER MET6 ;
        RECT 0 28.5 20 31.5 ;
      LAYER METG1 ;
        RECT 0 28.5 20 31.5 ;
      LAYER METS1 ;
        RECT 0 28.5 20 31.5 ;
      LAYER METS2 ;
        RECT 0 28.5 20 31.5 ;
      LAYER METS3 ;
        RECT 0 28.5 20 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 20 35.5 ;
      LAYER MET6 ;
        RECT 0 32.5 20 35.5 ;
      LAYER METG1 ;
        RECT 0 32.5 20 35.5 ;
      LAYER METS1 ;
        RECT 0 32.5 20 35.5 ;
      LAYER METS2 ;
        RECT 0 32.5 20 35.5 ;
      LAYER METS3 ;
        RECT 0 32.5 20 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 20 43.5 ;
      LAYER MET6 ;
        RECT 0 40.5 20 43.5 ;
      LAYER METG1 ;
        RECT 0 40.5 20 43.5 ;
      LAYER METS1 ;
        RECT 0 40.5 20 43.5 ;
      LAYER METS2 ;
        RECT 0 40.5 20 43.5 ;
      LAYER METS3 ;
        RECT 0 40.5 20 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 20 51.5 ;
      LAYER MET6 ;
        RECT 0 48.5 20 51.5 ;
      LAYER METG1 ;
        RECT 0 48.5 20 51.5 ;
      LAYER METS1 ;
        RECT 0 48.5 20 51.5 ;
      LAYER METS2 ;
        RECT 0 48.5 20 51.5 ;
      LAYER METS3 ;
        RECT 0 48.5 20 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 20 59.5 ;
      LAYER MET6 ;
        RECT 0 56.5 20 59.5 ;
      LAYER METG1 ;
        RECT 0 56.5 20 59.5 ;
      LAYER METS1 ;
        RECT 0 56.5 20 59.5 ;
      LAYER METS2 ;
        RECT 0 56.5 20 59.5 ;
      LAYER METS3 ;
        RECT 0 56.5 20 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 20 67.5 ;
      LAYER MET6 ;
        RECT 0 64.5 20 67.5 ;
      LAYER METG1 ;
        RECT 0 64.5 20 67.5 ;
      LAYER METS1 ;
        RECT 0 64.5 20 67.5 ;
      LAYER METS2 ;
        RECT 0 64.5 20 67.5 ;
      LAYER METS3 ;
        RECT 0 64.5 20 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 20 75.5 ;
      LAYER MET6 ;
        RECT 0 72.5 20 75.5 ;
      LAYER METG1 ;
        RECT 0 72.5 20 75.5 ;
      LAYER METS1 ;
        RECT 0 72.5 20 75.5 ;
      LAYER METS2 ;
        RECT 0 72.5 20 75.5 ;
      LAYER METS3 ;
        RECT 0 72.5 20 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 20 111.5 ;
      LAYER MET6 ;
        RECT 0 108.5 20 111.5 ;
      LAYER METG1 ;
        RECT 0 108.5 20 111.5 ;
      LAYER METS1 ;
        RECT 0 108.5 20 111.5 ;
      LAYER METS2 ;
        RECT 0 108.5 20 111.5 ;
      LAYER METS3 ;
        RECT 0 108.5 20 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 20 131.5 ;
      LAYER MET6 ;
        RECT 0 128.5 20 131.5 ;
      LAYER METG1 ;
        RECT 0 128.5 20 131.5 ;
      LAYER METS1 ;
        RECT 0 128.5 20 131.5 ;
      LAYER METS2 ;
        RECT 0 128.5 20 131.5 ;
      LAYER METS3 ;
        RECT 0 128.5 20 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 20 139.5 ;
      LAYER MET6 ;
        RECT 0 136.5 20 139.5 ;
      LAYER METG1 ;
        RECT 0 136.5 20 139.5 ;
      LAYER METS1 ;
        RECT 0 136.5 20 139.5 ;
      LAYER METS2 ;
        RECT 0 136.5 20 139.5 ;
      LAYER METS3 ;
        RECT 0 136.5 20 139.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 75.6 20 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 20 79.5 ;
      LAYER MET6 ;
        RECT 0 76.5 20 79.5 ;
      LAYER METG1 ;
        RECT 0 76.5 20 79.5 ;
      LAYER METS1 ;
        RECT 0 76.5 20 79.5 ;
      LAYER METS2 ;
        RECT 0 76.5 20 79.5 ;
      LAYER METS3 ;
        RECT 0 76.5 20 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 20 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 20 83.5 ;
      LAYER MET6 ;
        RECT 0 80.5 20 83.5 ;
      LAYER METG1 ;
        RECT 0 80.5 20 83.5 ;
      LAYER METS1 ;
        RECT 0 80.5 20 83.5 ;
      LAYER METS2 ;
        RECT 0 80.5 20 83.5 ;
      LAYER METS3 ;
        RECT 0 80.5 20 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 20 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 20 87.5 ;
      LAYER MET6 ;
        RECT 0 84.5 20 87.5 ;
      LAYER METG1 ;
        RECT 0 84.5 20 87.5 ;
      LAYER METS1 ;
        RECT 0 84.5 20 87.5 ;
      LAYER METS2 ;
        RECT 0 84.5 20 87.5 ;
      LAYER METS3 ;
        RECT 0 84.5 20 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 20 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 20 91.5 ;
      LAYER MET6 ;
        RECT 0 88.5 20 91.5 ;
      LAYER METG1 ;
        RECT 0 88.5 20 91.5 ;
      LAYER METS1 ;
        RECT 0 88.5 20 91.5 ;
      LAYER METS2 ;
        RECT 0 88.5 20 91.5 ;
      LAYER METS3 ;
        RECT 0 88.5 20 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 20 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 20 95.5 ;
      LAYER MET6 ;
        RECT 0 92.5 20 95.5 ;
      LAYER METG1 ;
        RECT 0 92.5 20 95.5 ;
      LAYER METS1 ;
        RECT 0 92.5 20 95.5 ;
      LAYER METS2 ;
        RECT 0 92.5 20 95.5 ;
      LAYER METS3 ;
        RECT 0 92.5 20 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 20 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 20 99.5 ;
      LAYER MET6 ;
        RECT 0 96.5 20 99.5 ;
      LAYER METG1 ;
        RECT 0 96.5 20 99.5 ;
      LAYER METS1 ;
        RECT 0 96.5 20 99.5 ;
      LAYER METS2 ;
        RECT 0 96.5 20 99.5 ;
      LAYER METS3 ;
        RECT 0 96.5 20 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 20 155.5 ;
      LAYER MET6 ;
        RECT 0 152.5 20 155.5 ;
      LAYER METG1 ;
        RECT 0 152.5 20 155.5 ;
      LAYER METS1 ;
        RECT 0 152.5 20 155.5 ;
      LAYER METS2 ;
        RECT 0 152.5 20 155.5 ;
      LAYER METS3 ;
        RECT 0 152.5 20 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 20 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 20 159.5 ;
      LAYER MET6 ;
        RECT 0 156.5 20 159.5 ;
      LAYER METG1 ;
        RECT 0 156.5 20 159.5 ;
      LAYER METS1 ;
        RECT 0 156.5 20 159.5 ;
      LAYER METS2 ;
        RECT 0 156.5 20 159.5 ;
      LAYER METS3 ;
        RECT 0 156.5 20 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 20 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 20 163.5 ;
      LAYER MET6 ;
        RECT 0 160.5 20 163.5 ;
      LAYER METG1 ;
        RECT 0 160.5 20 163.5 ;
      LAYER METS1 ;
        RECT 0 160.5 20 163.5 ;
      LAYER METS2 ;
        RECT 0 160.5 20 163.5 ;
      LAYER METS3 ;
        RECT 0 160.5 20 163.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 4.5 20 7.5 ;
      LAYER MET6 ;
        RECT 0 4.5 20 7.5 ;
      LAYER METG1 ;
        RECT 0 4.5 20 7.5 ;
      LAYER METS1 ;
        RECT 0 4.5 20 7.5 ;
      LAYER METS2 ;
        RECT 0 4.5 20 7.5 ;
      LAYER METS3 ;
        RECT 0 4.5 20 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 20 11.5 ;
      LAYER MET6 ;
        RECT 0 8.5 20 11.5 ;
      LAYER METG1 ;
        RECT 0 8.5 20 11.5 ;
      LAYER METS1 ;
        RECT 0 8.5 20 11.5 ;
      LAYER METS2 ;
        RECT 0 8.5 20 11.5 ;
      LAYER METS3 ;
        RECT 0 8.5 20 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 20 23.5 ;
      LAYER MET6 ;
        RECT 0 20.5 20 23.5 ;
      LAYER METG1 ;
        RECT 0 20.5 20 23.5 ;
      LAYER METS1 ;
        RECT 0 20.5 20 23.5 ;
      LAYER METS2 ;
        RECT 0 20.5 20 23.5 ;
      LAYER METS3 ;
        RECT 0 20.5 20 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 20 27.5 ;
      LAYER MET6 ;
        RECT 0 24.5 20 27.5 ;
      LAYER METG1 ;
        RECT 0 24.5 20 27.5 ;
      LAYER METS1 ;
        RECT 0 24.5 20 27.5 ;
      LAYER METS2 ;
        RECT 0 24.5 20 27.5 ;
      LAYER METS3 ;
        RECT 0 24.5 20 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 20 39.5 ;
      LAYER MET6 ;
        RECT 0 36.5 20 39.5 ;
      LAYER METG1 ;
        RECT 0 36.5 20 39.5 ;
      LAYER METS1 ;
        RECT 0 36.5 20 39.5 ;
      LAYER METS2 ;
        RECT 0 36.5 20 39.5 ;
      LAYER METS3 ;
        RECT 0 36.5 20 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 20 47.5 ;
      LAYER MET6 ;
        RECT 0 44.5 20 47.5 ;
      LAYER METG1 ;
        RECT 0 44.5 20 47.5 ;
      LAYER METS1 ;
        RECT 0 44.5 20 47.5 ;
      LAYER METS2 ;
        RECT 0 44.5 20 47.5 ;
      LAYER METS3 ;
        RECT 0 44.5 20 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 20 55.5 ;
      LAYER MET6 ;
        RECT 0 52.5 20 55.5 ;
      LAYER METG1 ;
        RECT 0 52.5 20 55.5 ;
      LAYER METS1 ;
        RECT 0 52.5 20 55.5 ;
      LAYER METS2 ;
        RECT 0 52.5 20 55.5 ;
      LAYER METS3 ;
        RECT 0 52.5 20 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 20 63.5 ;
      LAYER MET6 ;
        RECT 0 60.5 20 63.5 ;
      LAYER METG1 ;
        RECT 0 60.5 20 63.5 ;
      LAYER METS1 ;
        RECT 0 60.5 20 63.5 ;
      LAYER METS2 ;
        RECT 0 60.5 20 63.5 ;
      LAYER METS3 ;
        RECT 0 60.5 20 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 20 71.5 ;
      LAYER MET6 ;
        RECT 0 68.5 20 71.5 ;
      LAYER METG1 ;
        RECT 0 68.5 20 71.5 ;
      LAYER METS1 ;
        RECT 0 68.5 20 71.5 ;
      LAYER METS2 ;
        RECT 0 68.5 20 71.5 ;
      LAYER METS3 ;
        RECT 0 68.5 20 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 20 103.5 ;
      LAYER MET6 ;
        RECT 0 100.5 20 103.5 ;
      LAYER METG1 ;
        RECT 0 100.5 20 103.5 ;
      LAYER METS1 ;
        RECT 0 100.5 20 103.5 ;
      LAYER METS2 ;
        RECT 0 100.5 20 103.5 ;
      LAYER METS3 ;
        RECT 0 100.5 20 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 20 135.5 ;
      LAYER MET6 ;
        RECT 0 132.5 20 135.5 ;
      LAYER METG1 ;
        RECT 0 132.5 20 135.5 ;
      LAYER METS1 ;
        RECT 0 132.5 20 135.5 ;
      LAYER METS2 ;
        RECT 0 132.5 20 135.5 ;
      LAYER METS3 ;
        RECT 0 132.5 20 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 103.6 20 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 20 107.5 ;
      LAYER MET6 ;
        RECT 0 104.5 20 107.5 ;
      LAYER METG1 ;
        RECT 0 104.5 20 107.5 ;
      LAYER METS1 ;
        RECT 0 104.5 20 107.5 ;
      LAYER METS2 ;
        RECT 0 104.5 20 107.5 ;
      LAYER METS3 ;
        RECT 0 104.5 20 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 20 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 20 115.5 ;
      LAYER MET6 ;
        RECT 0 112.5 20 115.5 ;
      LAYER METG1 ;
        RECT 0 112.5 20 115.5 ;
      LAYER METS1 ;
        RECT 0 112.5 20 115.5 ;
      LAYER METS2 ;
        RECT 0 112.5 20 115.5 ;
      LAYER METS3 ;
        RECT 0 112.5 20 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 20 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 20 119.5 ;
      LAYER MET6 ;
        RECT 0 116.5 20 119.5 ;
      LAYER METG1 ;
        RECT 0 116.5 20 119.5 ;
      LAYER METS1 ;
        RECT 0 116.5 20 119.5 ;
      LAYER METS2 ;
        RECT 0 116.5 20 119.5 ;
      LAYER METS3 ;
        RECT 0 116.5 20 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 20 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 20 123.5 ;
      LAYER MET6 ;
        RECT 0 120.5 20 123.5 ;
      LAYER METG1 ;
        RECT 0 120.5 20 123.5 ;
      LAYER METS1 ;
        RECT 0 120.5 20 123.5 ;
      LAYER METS2 ;
        RECT 0 120.5 20 123.5 ;
      LAYER METS3 ;
        RECT 0 120.5 20 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 20 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 20 127.5 ;
      LAYER MET6 ;
        RECT 0 124.5 20 127.5 ;
      LAYER METG1 ;
        RECT 0 124.5 20 127.5 ;
      LAYER METS1 ;
        RECT 0 124.5 20 127.5 ;
      LAYER METS2 ;
        RECT 0 124.5 20 127.5 ;
      LAYER METS3 ;
        RECT 0 124.5 20 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 20 143.5 ;
      LAYER MET6 ;
        RECT 0 140.5 20 143.5 ;
      LAYER METG1 ;
        RECT 0 140.5 20 143.5 ;
      LAYER METS1 ;
        RECT 0 140.5 20 143.5 ;
      LAYER METS2 ;
        RECT 0 140.5 20 143.5 ;
      LAYER METS3 ;
        RECT 0 140.5 20 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 20 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 20 147.5 ;
      LAYER MET6 ;
        RECT 0 144.5 20 147.5 ;
      LAYER METG1 ;
        RECT 0 144.5 20 147.5 ;
      LAYER METS1 ;
        RECT 0 144.5 20 147.5 ;
      LAYER METS2 ;
        RECT 0 144.5 20 147.5 ;
      LAYER METS3 ;
        RECT 0 144.5 20 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 20 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 20 151.5 ;
      LAYER MET6 ;
        RECT 0 148.5 20 151.5 ;
      LAYER METG1 ;
        RECT 0 148.5 20 151.5 ;
      LAYER METS1 ;
        RECT 0 148.5 20 151.5 ;
      LAYER METS2 ;
        RECT 0 148.5 20 151.5 ;
      LAYER METS3 ;
        RECT 0 148.5 20 151.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 20 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 20 15.5 ;
      LAYER MET6 ;
        RECT 0 12.5 20 15.5 ;
      LAYER METG1 ;
        RECT 0 12.5 20 15.5 ;
      LAYER METS1 ;
        RECT 0 12.5 20 15.5 ;
      LAYER METS2 ;
        RECT 0 12.5 20 15.5 ;
      LAYER METS3 ;
        RECT 0 12.5 20 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 20 19.5 ;
      LAYER MET6 ;
        RECT 0 16.5 20 19.5 ;
      LAYER METG1 ;
        RECT 0 16.5 20 19.5 ;
      LAYER METS1 ;
        RECT 0 16.5 20 19.5 ;
      LAYER METS2 ;
        RECT 0 16.5 20 19.5 ;
      LAYER METS3 ;
        RECT 0 16.5 20 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 20 170 ;
    LAYER CUT12 ;
      RECT 0 0 20 170 ;
    LAYER MET2 ;
      RECT 0 0 20 170 ;
    LAYER CUT23 ;
      RECT 0 0 20 170 ;
    LAYER MET3 ;
      RECT 0 0 20 170 ;
    LAYER CUT34 ;
      RECT 0 0 20 170 ;
    LAYER MET4 ;
      RECT 0 0 20 170 ;
    LAYER CUT45 ;
      RECT 0 0 20 170 ;
    LAYER MET5 ;
      RECT 0 0 20 170 ;
    LAYER CUT56 ;
      RECT 0 0 20 170 ;
    LAYER MET6 ;
      RECT 0 0 20 170 ;
    LAYER CUTS1 ;
      RECT 0 0 20 170 ;
    LAYER METS1 ;
      RECT 0 0 20 170 ;
    LAYER CUTS2 ;
      RECT 0 0 20 170 ;
    LAYER METS2 ;
      RECT 0 0 20 170 ;
    LAYER CUTS3 ;
      RECT 0 0 20 170 ;
    LAYER METS3 ;
      RECT 0 0 20 170 ;
    LAYER CUTG1 ;
      RECT 0 0 20 170 ;
    LAYER METG1 ;
      RECT 0 0 20 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 20.000 2.000 ;
  END
END IOCB2ESD4C0A1


MACRO IOCB2ESE4C0A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2ESE4C0A1 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 28.5 40 31.5 ;
      LAYER MET6 ;
        RECT 0 28.5 40 31.5 ;
      LAYER METG1 ;
        RECT 0 28.5 40 31.5 ;
      LAYER METS1 ;
        RECT 0 28.5 40 31.5 ;
      LAYER METS2 ;
        RECT 0 28.5 40 31.5 ;
      LAYER METS3 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 32.5 40 35.5 ;
      LAYER MET6 ;
        RECT 0 32.5 40 35.5 ;
      LAYER METG1 ;
        RECT 0 32.5 40 35.5 ;
      LAYER METS1 ;
        RECT 0 32.5 40 35.5 ;
      LAYER METS2 ;
        RECT 0 32.5 40 35.5 ;
      LAYER METS3 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 40.5 40 43.5 ;
      LAYER MET6 ;
        RECT 0 40.5 40 43.5 ;
      LAYER METG1 ;
        RECT 0 40.5 40 43.5 ;
      LAYER METS1 ;
        RECT 0 40.5 40 43.5 ;
      LAYER METS2 ;
        RECT 0 40.5 40 43.5 ;
      LAYER METS3 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 48.5 40 51.5 ;
      LAYER MET6 ;
        RECT 0 48.5 40 51.5 ;
      LAYER METG1 ;
        RECT 0 48.5 40 51.5 ;
      LAYER METS1 ;
        RECT 0 48.5 40 51.5 ;
      LAYER METS2 ;
        RECT 0 48.5 40 51.5 ;
      LAYER METS3 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 56.5 40 59.5 ;
      LAYER MET6 ;
        RECT 0 56.5 40 59.5 ;
      LAYER METG1 ;
        RECT 0 56.5 40 59.5 ;
      LAYER METS1 ;
        RECT 0 56.5 40 59.5 ;
      LAYER METS2 ;
        RECT 0 56.5 40 59.5 ;
      LAYER METS3 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 64.5 40 67.5 ;
      LAYER MET6 ;
        RECT 0 64.5 40 67.5 ;
      LAYER METG1 ;
        RECT 0 64.5 40 67.5 ;
      LAYER METS1 ;
        RECT 0 64.5 40 67.5 ;
      LAYER METS2 ;
        RECT 0 64.5 40 67.5 ;
      LAYER METS3 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 72.5 40 75.5 ;
      LAYER MET6 ;
        RECT 0 72.5 40 75.5 ;
      LAYER METG1 ;
        RECT 0 72.5 40 75.5 ;
      LAYER METS1 ;
        RECT 0 72.5 40 75.5 ;
      LAYER METS2 ;
        RECT 0 72.5 40 75.5 ;
      LAYER METS3 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 108.5 40 111.5 ;
      LAYER MET6 ;
        RECT 0 108.5 40 111.5 ;
      LAYER METG1 ;
        RECT 0 108.5 40 111.5 ;
      LAYER METS1 ;
        RECT 0 108.5 40 111.5 ;
      LAYER METS2 ;
        RECT 0 108.5 40 111.5 ;
      LAYER METS3 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 128.5 40 131.5 ;
      LAYER MET6 ;
        RECT 0 128.5 40 131.5 ;
      LAYER METG1 ;
        RECT 0 128.5 40 131.5 ;
      LAYER METS1 ;
        RECT 0 128.5 40 131.5 ;
      LAYER METS2 ;
        RECT 0 128.5 40 131.5 ;
      LAYER METS3 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 136.5 40 139.5 ;
      LAYER MET6 ;
        RECT 0 136.5 40 139.5 ;
      LAYER METG1 ;
        RECT 0 136.5 40 139.5 ;
      LAYER METS1 ;
        RECT 0 136.5 40 139.5 ;
      LAYER METS2 ;
        RECT 0 136.5 40 139.5 ;
      LAYER METS3 ;
        RECT 0 136.5 40 139.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 75.6 40 78.6 ;
      LAYER MET5 ;
        RECT 0 76.5 40 79.5 ;
      LAYER MET6 ;
        RECT 0 76.5 40 79.5 ;
      LAYER METG1 ;
        RECT 0 76.5 40 79.5 ;
      LAYER METS1 ;
        RECT 0 76.5 40 79.5 ;
      LAYER METS2 ;
        RECT 0 76.5 40 79.5 ;
      LAYER METS3 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 79.6 40 82.6 ;
      LAYER MET5 ;
        RECT 0 80.5 40 83.5 ;
      LAYER MET6 ;
        RECT 0 80.5 40 83.5 ;
      LAYER METG1 ;
        RECT 0 80.5 40 83.5 ;
      LAYER METS1 ;
        RECT 0 80.5 40 83.5 ;
      LAYER METS2 ;
        RECT 0 80.5 40 83.5 ;
      LAYER METS3 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 83.6 40 86.6 ;
      LAYER MET5 ;
        RECT 0 84.5 40 87.5 ;
      LAYER MET6 ;
        RECT 0 84.5 40 87.5 ;
      LAYER METG1 ;
        RECT 0 84.5 40 87.5 ;
      LAYER METS1 ;
        RECT 0 84.5 40 87.5 ;
      LAYER METS2 ;
        RECT 0 84.5 40 87.5 ;
      LAYER METS3 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 87.6 40 90.6 ;
      LAYER MET5 ;
        RECT 0 88.5 40 91.5 ;
      LAYER MET6 ;
        RECT 0 88.5 40 91.5 ;
      LAYER METG1 ;
        RECT 0 88.5 40 91.5 ;
      LAYER METS1 ;
        RECT 0 88.5 40 91.5 ;
      LAYER METS2 ;
        RECT 0 88.5 40 91.5 ;
      LAYER METS3 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 91.6 40 94.6 ;
      LAYER MET5 ;
        RECT 0 92.5 40 95.5 ;
      LAYER MET6 ;
        RECT 0 92.5 40 95.5 ;
      LAYER METG1 ;
        RECT 0 92.5 40 95.5 ;
      LAYER METS1 ;
        RECT 0 92.5 40 95.5 ;
      LAYER METS2 ;
        RECT 0 92.5 40 95.5 ;
      LAYER METS3 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 95.6 40 98.6 ;
      LAYER MET5 ;
        RECT 0 96.5 40 99.5 ;
      LAYER MET6 ;
        RECT 0 96.5 40 99.5 ;
      LAYER METG1 ;
        RECT 0 96.5 40 99.5 ;
      LAYER METS1 ;
        RECT 0 96.5 40 99.5 ;
      LAYER METS2 ;
        RECT 0 96.5 40 99.5 ;
      LAYER METS3 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET6 ;
        RECT 0 152.5 40 155.5 ;
      LAYER METG1 ;
        RECT 0 152.5 40 155.5 ;
      LAYER METS1 ;
        RECT 0 152.5 40 155.5 ;
      LAYER METS2 ;
        RECT 0 152.5 40 155.5 ;
      LAYER METS3 ;
        RECT 0 152.5 40 155.5 ;
      LAYER MET3 ;
        RECT 0 153.43 40 156.43 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET6 ;
        RECT 0 156.5 40 159.5 ;
      LAYER METG1 ;
        RECT 0 156.5 40 159.5 ;
      LAYER METS1 ;
        RECT 0 156.5 40 159.5 ;
      LAYER METS2 ;
        RECT 0 156.5 40 159.5 ;
      LAYER METS3 ;
        RECT 0 156.5 40 159.5 ;
      LAYER MET3 ;
        RECT 0 158.99 40 161.99 ;
      LAYER MET5 ;
        RECT 0 160.5 40 163.5 ;
      LAYER MET6 ;
        RECT 0 160.5 40 163.5 ;
      LAYER METG1 ;
        RECT 0 160.5 40 163.5 ;
      LAYER METS1 ;
        RECT 0 160.5 40 163.5 ;
      LAYER METS2 ;
        RECT 0 160.5 40 163.5 ;
      LAYER METS3 ;
        RECT 0 160.5 40 163.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 4.5 40 7.5 ;
      LAYER MET6 ;
        RECT 0 4.5 40 7.5 ;
      LAYER METG1 ;
        RECT 0 4.5 40 7.5 ;
      LAYER METS1 ;
        RECT 0 4.5 40 7.5 ;
      LAYER METS2 ;
        RECT 0 4.5 40 7.5 ;
      LAYER METS3 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 8.5 40 11.5 ;
      LAYER MET6 ;
        RECT 0 8.5 40 11.5 ;
      LAYER METG1 ;
        RECT 0 8.5 40 11.5 ;
      LAYER METS1 ;
        RECT 0 8.5 40 11.5 ;
      LAYER METS2 ;
        RECT 0 8.5 40 11.5 ;
      LAYER METS3 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 20.5 40 23.5 ;
      LAYER MET6 ;
        RECT 0 20.5 40 23.5 ;
      LAYER METG1 ;
        RECT 0 20.5 40 23.5 ;
      LAYER METS1 ;
        RECT 0 20.5 40 23.5 ;
      LAYER METS2 ;
        RECT 0 20.5 40 23.5 ;
      LAYER METS3 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 24.5 40 27.5 ;
      LAYER MET6 ;
        RECT 0 24.5 40 27.5 ;
      LAYER METG1 ;
        RECT 0 24.5 40 27.5 ;
      LAYER METS1 ;
        RECT 0 24.5 40 27.5 ;
      LAYER METS2 ;
        RECT 0 24.5 40 27.5 ;
      LAYER METS3 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 36.5 40 39.5 ;
      LAYER MET6 ;
        RECT 0 36.5 40 39.5 ;
      LAYER METG1 ;
        RECT 0 36.5 40 39.5 ;
      LAYER METS1 ;
        RECT 0 36.5 40 39.5 ;
      LAYER METS2 ;
        RECT 0 36.5 40 39.5 ;
      LAYER METS3 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 44.5 40 47.5 ;
      LAYER MET6 ;
        RECT 0 44.5 40 47.5 ;
      LAYER METG1 ;
        RECT 0 44.5 40 47.5 ;
      LAYER METS1 ;
        RECT 0 44.5 40 47.5 ;
      LAYER METS2 ;
        RECT 0 44.5 40 47.5 ;
      LAYER METS3 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 52.5 40 55.5 ;
      LAYER MET6 ;
        RECT 0 52.5 40 55.5 ;
      LAYER METG1 ;
        RECT 0 52.5 40 55.5 ;
      LAYER METS1 ;
        RECT 0 52.5 40 55.5 ;
      LAYER METS2 ;
        RECT 0 52.5 40 55.5 ;
      LAYER METS3 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 60.5 40 63.5 ;
      LAYER MET6 ;
        RECT 0 60.5 40 63.5 ;
      LAYER METG1 ;
        RECT 0 60.5 40 63.5 ;
      LAYER METS1 ;
        RECT 0 60.5 40 63.5 ;
      LAYER METS2 ;
        RECT 0 60.5 40 63.5 ;
      LAYER METS3 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 68.5 40 71.5 ;
      LAYER MET6 ;
        RECT 0 68.5 40 71.5 ;
      LAYER METG1 ;
        RECT 0 68.5 40 71.5 ;
      LAYER METS1 ;
        RECT 0 68.5 40 71.5 ;
      LAYER METS2 ;
        RECT 0 68.5 40 71.5 ;
      LAYER METS3 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 100.5 40 103.5 ;
      LAYER MET6 ;
        RECT 0 100.5 40 103.5 ;
      LAYER METG1 ;
        RECT 0 100.5 40 103.5 ;
      LAYER METS1 ;
        RECT 0 100.5 40 103.5 ;
      LAYER METS2 ;
        RECT 0 100.5 40 103.5 ;
      LAYER METS3 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 132.5 40 135.5 ;
      LAYER MET6 ;
        RECT 0 132.5 40 135.5 ;
      LAYER METG1 ;
        RECT 0 132.5 40 135.5 ;
      LAYER METS1 ;
        RECT 0 132.5 40 135.5 ;
      LAYER METS2 ;
        RECT 0 132.5 40 135.5 ;
      LAYER METS3 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 103.6 40 106.6 ;
      LAYER MET5 ;
        RECT 0 104.5 40 107.5 ;
      LAYER MET6 ;
        RECT 0 104.5 40 107.5 ;
      LAYER METG1 ;
        RECT 0 104.5 40 107.5 ;
      LAYER METS1 ;
        RECT 0 104.5 40 107.5 ;
      LAYER METS2 ;
        RECT 0 104.5 40 107.5 ;
      LAYER METS3 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 111.6 40 114.6 ;
      LAYER MET5 ;
        RECT 0 112.5 40 115.5 ;
      LAYER MET6 ;
        RECT 0 112.5 40 115.5 ;
      LAYER METG1 ;
        RECT 0 112.5 40 115.5 ;
      LAYER METS1 ;
        RECT 0 112.5 40 115.5 ;
      LAYER METS2 ;
        RECT 0 112.5 40 115.5 ;
      LAYER METS3 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 115.6 40 118.6 ;
      LAYER MET5 ;
        RECT 0 116.5 40 119.5 ;
      LAYER MET6 ;
        RECT 0 116.5 40 119.5 ;
      LAYER METG1 ;
        RECT 0 116.5 40 119.5 ;
      LAYER METS1 ;
        RECT 0 116.5 40 119.5 ;
      LAYER METS2 ;
        RECT 0 116.5 40 119.5 ;
      LAYER METS3 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 119.6 40 122.6 ;
      LAYER MET5 ;
        RECT 0 120.5 40 123.5 ;
      LAYER MET6 ;
        RECT 0 120.5 40 123.5 ;
      LAYER METG1 ;
        RECT 0 120.5 40 123.5 ;
      LAYER METS1 ;
        RECT 0 120.5 40 123.5 ;
      LAYER METS2 ;
        RECT 0 120.5 40 123.5 ;
      LAYER METS3 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 123.6 40 126.6 ;
      LAYER MET5 ;
        RECT 0 124.5 40 127.5 ;
      LAYER MET6 ;
        RECT 0 124.5 40 127.5 ;
      LAYER METG1 ;
        RECT 0 124.5 40 127.5 ;
      LAYER METS1 ;
        RECT 0 124.5 40 127.5 ;
      LAYER METS2 ;
        RECT 0 124.5 40 127.5 ;
      LAYER METS3 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET6 ;
        RECT 0 140.5 40 143.5 ;
      LAYER METG1 ;
        RECT 0 140.5 40 143.5 ;
      LAYER METS1 ;
        RECT 0 140.5 40 143.5 ;
      LAYER METS2 ;
        RECT 0 140.5 40 143.5 ;
      LAYER METS3 ;
        RECT 0 140.5 40 143.5 ;
      LAYER MET3 ;
        RECT 0 142.84 40 145.84 ;
      LAYER MET5 ;
        RECT 0 144.5 40 147.5 ;
      LAYER MET6 ;
        RECT 0 144.5 40 147.5 ;
      LAYER METG1 ;
        RECT 0 144.5 40 147.5 ;
      LAYER METS1 ;
        RECT 0 144.5 40 147.5 ;
      LAYER METS2 ;
        RECT 0 144.5 40 147.5 ;
      LAYER METS3 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 148.4 40 151.4 ;
      LAYER MET5 ;
        RECT 0 148.5 40 151.5 ;
      LAYER MET6 ;
        RECT 0 148.5 40 151.5 ;
      LAYER METG1 ;
        RECT 0 148.5 40 151.5 ;
      LAYER METS1 ;
        RECT 0 148.5 40 151.5 ;
      LAYER METS2 ;
        RECT 0 148.5 40 151.5 ;
      LAYER METS3 ;
        RECT 0 148.5 40 151.5 ;
    END
    PORT
      LAYER MET3 ;
        RECT 0 107.6 40 110.6 ;
    END
  END VSS
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET5 ;
        RECT 0 12.5 40 15.5 ;
      LAYER MET6 ;
        RECT 0 12.5 40 15.5 ;
      LAYER METG1 ;
        RECT 0 12.5 40 15.5 ;
      LAYER METS1 ;
        RECT 0 12.5 40 15.5 ;
      LAYER METS2 ;
        RECT 0 12.5 40 15.5 ;
      LAYER METS3 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET5 ;
        RECT 0 16.5 40 19.5 ;
      LAYER MET6 ;
        RECT 0 16.5 40 19.5 ;
      LAYER METG1 ;
        RECT 0 16.5 40 19.5 ;
      LAYER METS1 ;
        RECT 0 16.5 40 19.5 ;
      LAYER METS2 ;
        RECT 0 16.5 40 19.5 ;
      LAYER METS3 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  OBS
    LAYER MET1 ;
      RECT 0 0 40 170 ;
    LAYER CUT12 ;
      RECT 0 0 40 170 ;
    LAYER MET2 ;
      RECT 0 0 40 170 ;
    LAYER CUT23 ;
      RECT 0 0 40 170 ;
    LAYER MET3 ;
      RECT 0 0 40 170 ;
    LAYER CUT34 ;
      RECT 0 0 40 170 ;
    LAYER MET4 ;
      RECT 0 0 40 170 ;
    LAYER CUT45 ;
      RECT 0 0 40 170 ;
    LAYER MET5 ;
      RECT 0 0 40 170 ;
    LAYER CUT56 ;
      RECT 0 0 40 170 ;
    LAYER MET6 ;
      RECT 0 0 40 170 ;
    LAYER CUTS1 ;
      RECT 0 0 40 170 ;
    LAYER METS1 ;
      RECT 0 0 40 170 ;
    LAYER CUTS2 ;
      RECT 0 0 40 170 ;
    LAYER METS2 ;
      RECT 0 0 40 170 ;
    LAYER CUTS3 ;
      RECT 0 0 40 170 ;
    LAYER METS3 ;
      RECT 0 0 40 170 ;
    LAYER CUTG1 ;
      RECT 0 0 40 170 ;
    LAYER METG1 ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 0.000 40.000 2.000 ;
  END
END IOCB2ESE4C0A1


MACRO IOCB2EW3A5C0A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EW3A5C0A1 0 0 ;
  SIZE 50 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET6 ;
        RECT 0 12.5 50 15.5 ;
      LAYER METG1 ;
        RECT 0 12.5 50 15.5 ;
      LAYER METS2 ;
        RECT 0 12.5 50 15.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 16.5 50 19.5 ;
      LAYER METG1 ;
        RECT 0 16.5 50 19.5 ;
      LAYER METS2 ;
        RECT 0 16.5 50 19.5 ;
    END
  END VDD
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET6 ;
        RECT 0 28.5 50 31.5 ;
      LAYER METG1 ;
        RECT 0 28.5 50 31.5 ;
      LAYER METS2 ;
        RECT 0 28.5 50 31.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 32.5 50 35.5 ;
      LAYER METG1 ;
        RECT 0 32.5 50 35.5 ;
      LAYER METS2 ;
        RECT 0 32.5 50 35.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 40.5 50 43.5 ;
      LAYER METG1 ;
        RECT 0 40.5 50 43.5 ;
      LAYER METS2 ;
        RECT 0 40.5 50 43.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 48.5 50 51.5 ;
      LAYER METG1 ;
        RECT 0 48.5 50 51.5 ;
      LAYER METS2 ;
        RECT 0 48.5 50 51.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 56.5 50 59.5 ;
      LAYER METG1 ;
        RECT 0 56.5 50 59.5 ;
      LAYER METS2 ;
        RECT 0 56.5 50 59.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 64.5 50 67.5 ;
      LAYER METG1 ;
        RECT 0 64.5 50 67.5 ;
      LAYER METS2 ;
        RECT 0 64.5 50 67.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 72.5 50 75.5 ;
      LAYER METG1 ;
        RECT 0 72.5 50 75.5 ;
      LAYER METS2 ;
        RECT 0 72.5 50 75.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 76.5 50 79.5 ;
      LAYER METG1 ;
        RECT 0 76.5 50 79.5 ;
      LAYER METS2 ;
        RECT 0 76.5 50 79.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 80.5 50 83.5 ;
      LAYER METG1 ;
        RECT 0 80.5 50 83.5 ;
      LAYER METS2 ;
        RECT 0 80.5 50 83.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 84.5 50 87.5 ;
      LAYER METG1 ;
        RECT 0 84.5 50 87.5 ;
      LAYER METS2 ;
        RECT 0 84.5 50 87.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 88.5 50 91.5 ;
      LAYER METG1 ;
        RECT 0 88.5 50 91.5 ;
      LAYER METS2 ;
        RECT 0 88.5 50 91.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 92.5 50 95.5 ;
      LAYER METG1 ;
        RECT 0 92.5 50 95.5 ;
      LAYER METS2 ;
        RECT 0 92.5 50 95.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 96.5 50 99.5 ;
      LAYER METG1 ;
        RECT 0 96.5 50 99.5 ;
      LAYER METS2 ;
        RECT 0 96.5 50 99.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 108.5 50 111.5 ;
      LAYER METG1 ;
        RECT 0 108.5 50 111.5 ;
      LAYER METS2 ;
        RECT 0 108.5 50 111.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 128.5 50 131.5 ;
      LAYER METG1 ;
        RECT 0 128.5 50 131.5 ;
      LAYER METS2 ;
        RECT 0 128.5 50 131.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 136.5 50 139.5 ;
      LAYER METG1 ;
        RECT 0 136.5 50 139.5 ;
      LAYER METS2 ;
        RECT 0 136.5 50 139.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 152.5 50 155.5 ;
      LAYER METG1 ;
        RECT 0 152.5 50 155.5 ;
      LAYER METS2 ;
        RECT 0 152.5 50 155.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 156.5 50 159.5 ;
      LAYER METG1 ;
        RECT 0 156.5 50 159.5 ;
      LAYER METS2 ;
        RECT 0 156.5 50 159.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 160.5 50 163.5 ;
      LAYER METG1 ;
        RECT 0 160.5 50 163.5 ;
      LAYER METS2 ;
        RECT 0 160.5 50 163.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET6 ;
        RECT 0 4.5 50 7.5 ;
      LAYER METG1 ;
        RECT 0 4.5 50 7.5 ;
      LAYER METS2 ;
        RECT 0 4.5 50 7.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 8.5 50 11.5 ;
      LAYER METG1 ;
        RECT 0 8.5 50 11.5 ;
      LAYER METS2 ;
        RECT 0 8.5 50 11.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 20.5 50 23.5 ;
      LAYER METG1 ;
        RECT 0 20.5 50 23.5 ;
      LAYER METS2 ;
        RECT 0 20.5 50 23.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 24.5 50 27.5 ;
      LAYER METG1 ;
        RECT 0 24.5 50 27.5 ;
      LAYER METS2 ;
        RECT 0 24.5 50 27.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 36.5 50 39.5 ;
      LAYER METG1 ;
        RECT 0 36.5 50 39.5 ;
      LAYER METS2 ;
        RECT 0 36.5 50 39.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 44.5 50 47.5 ;
      LAYER METG1 ;
        RECT 0 44.5 50 47.5 ;
      LAYER METS2 ;
        RECT 0 44.5 50 47.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 52.5 50 55.5 ;
      LAYER METG1 ;
        RECT 0 52.5 50 55.5 ;
      LAYER METS2 ;
        RECT 0 52.5 50 55.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 60.5 50 63.5 ;
      LAYER METG1 ;
        RECT 0 60.5 50 63.5 ;
      LAYER METS2 ;
        RECT 0 60.5 50 63.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 68.5 50 71.5 ;
      LAYER METG1 ;
        RECT 0 68.5 50 71.5 ;
      LAYER METS2 ;
        RECT 0 68.5 50 71.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 100.5 50 103.5 ;
      LAYER METG1 ;
        RECT 0 100.5 50 103.5 ;
      LAYER METS2 ;
        RECT 0 100.5 50 103.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 104.5 50 107.5 ;
      LAYER METG1 ;
        RECT 0 104.5 50 107.5 ;
      LAYER METS2 ;
        RECT 0 104.5 50 107.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 112.5 50 115.5 ;
      LAYER METG1 ;
        RECT 0 112.5 50 115.5 ;
      LAYER METS2 ;
        RECT 0 112.5 50 115.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 116.5 50 119.5 ;
      LAYER METG1 ;
        RECT 0 116.5 50 119.5 ;
      LAYER METS2 ;
        RECT 0 116.5 50 119.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 120.5 50 123.5 ;
      LAYER METG1 ;
        RECT 0 120.5 50 123.5 ;
      LAYER METS2 ;
        RECT 0 120.5 50 123.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 124.5 50 127.5 ;
      LAYER METG1 ;
        RECT 0 124.5 50 127.5 ;
      LAYER METS2 ;
        RECT 0 124.5 50 127.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 132.5 50 135.5 ;
      LAYER METG1 ;
        RECT 0 132.5 50 135.5 ;
      LAYER METS2 ;
        RECT 0 132.5 50 135.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 140.5 50 143.5 ;
      LAYER METG1 ;
        RECT 0 140.5 50 143.5 ;
      LAYER METS2 ;
        RECT 0 140.5 50 143.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 144.5 50 147.5 ;
      LAYER METG1 ;
        RECT 0 144.5 50 147.5 ;
      LAYER METS2 ;
        RECT 0 144.5 50 147.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 148.5 50 151.5 ;
      LAYER METG1 ;
        RECT 0 148.5 50 151.5 ;
      LAYER METS2 ;
        RECT 0 148.5 50 151.5 ;
    END
  END VSS
  OBS
    LAYER CUT56 ;
      RECT 0 0 50 170 ;
    LAYER MET6 ;
      RECT 0 0 50 170 ;
    LAYER CUTS1 ;
      RECT 0 0 50 170 ;
    LAYER METS1 ;
      RECT 0 0 50 170 ;
    LAYER CUTS2 ;
      RECT 0 0 50 170 ;
    LAYER METS2 ;
      RECT 0 0 50 170 ;
    LAYER CUTS3 ;
      RECT 0 0 50 170 ;
    LAYER METS3 ;
      RECT 0 0 50 170 ;
    LAYER CUTG1 ;
      RECT 0 0 50 170 ;
    LAYER METG1 ;
      RECT 0 0 50 170 ;
    LAYER CUTG2 ;
      RECT 0 0 50 170 ;
    LAYER METG2 ;
      RECT 0 0 50 170 ;
    LAYER CUTTOP ;
      RECT 0 0 50 170 ;
    LAYER METTOP ;
      RECT 0 0 50 170 ;
      LAYER OVLAP ;
       RECT 0.000 84.000 50.000 86.000 ;
  END
END IOCB2EW3A5C0A1


MACRO IOCB2EWDA5C0A1
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EWDA5C0A1 0 0 ;
  SIZE 50 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      CLASS CORE ;
      LAYER METG2 ;
        RECT 14.5 0 20.5 5 ;
      LAYER METTOP ;
        RECT 14.5 0 20.5 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG2 ;
        RECT 22 0 28 5 ;
      LAYER METTOP ;
        RECT 22 0 28 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG2 ;
        RECT 29.5 0 35.5 5 ;
      LAYER METTOP ;
        RECT 29.5 0 35.5 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG2 ;
        RECT 37 0 43 5 ;
      LAYER METTOP ;
        RECT 37 0 43 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG2 ;
        RECT 7 0 13 5 ;
      LAYER METTOP ;
        RECT 7 0 13 5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 12.5 50 15.5 ;
      LAYER METG1 ;
        RECT 0 12.5 50 15.5 ;
      LAYER METS2 ;
        RECT 0 12.5 50 15.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 16.5 50 19.5 ;
      LAYER METG1 ;
        RECT 0 16.5 50 19.5 ;
      LAYER METS2 ;
        RECT 0 16.5 50 19.5 ;
    END
  END VDD
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET6 ;
        RECT 0 28.5 50 31.5 ;
      LAYER METG1 ;
        RECT 0 28.5 50 31.5 ;
      LAYER METS2 ;
        RECT 0 28.5 50 31.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 32.5 50 35.5 ;
      LAYER METG1 ;
        RECT 0 32.5 50 35.5 ;
      LAYER METS2 ;
        RECT 0 32.5 50 35.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 40.5 50 43.5 ;
      LAYER METG1 ;
        RECT 0 40.5 50 43.5 ;
      LAYER METS2 ;
        RECT 0 40.5 50 43.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 48.5 50 51.5 ;
      LAYER METG1 ;
        RECT 0 48.5 50 51.5 ;
      LAYER METS2 ;
        RECT 0 48.5 50 51.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 56.5 50 59.5 ;
      LAYER METG1 ;
        RECT 0 56.5 50 59.5 ;
      LAYER METS2 ;
        RECT 0 56.5 50 59.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 64.5 50 67.5 ;
      LAYER METG1 ;
        RECT 0 64.5 50 67.5 ;
      LAYER METS2 ;
        RECT 0 64.5 50 67.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 72.5 50 75.5 ;
      LAYER METG1 ;
        RECT 0 72.5 50 75.5 ;
      LAYER METS2 ;
        RECT 0 72.5 50 75.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 76.5 50 79.5 ;
      LAYER METG1 ;
        RECT 0 76.5 50 79.5 ;
      LAYER METS2 ;
        RECT 0 76.5 50 79.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 80.5 50 83.5 ;
      LAYER METG1 ;
        RECT 0 80.5 50 83.5 ;
      LAYER METS2 ;
        RECT 0 80.5 50 83.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 84.5 50 87.5 ;
      LAYER METG1 ;
        RECT 0 84.5 50 87.5 ;
      LAYER METS2 ;
        RECT 0 84.5 50 87.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 88.5 50 91.5 ;
      LAYER METG1 ;
        RECT 0 88.5 50 91.5 ;
      LAYER METS2 ;
        RECT 0 88.5 50 91.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 92.5 50 95.5 ;
      LAYER METG1 ;
        RECT 0 92.5 50 95.5 ;
      LAYER METS2 ;
        RECT 0 92.5 50 95.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 96.5 50 99.5 ;
      LAYER METG1 ;
        RECT 0 96.5 50 99.5 ;
      LAYER METS2 ;
        RECT 0 96.5 50 99.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 108.5 50 111.5 ;
      LAYER METG1 ;
        RECT 0 108.5 50 111.5 ;
      LAYER METS2 ;
        RECT 0 108.5 50 111.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 128.5 50 131.5 ;
      LAYER METG1 ;
        RECT 0 128.5 50 131.5 ;
      LAYER METS2 ;
        RECT 0 128.5 50 131.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 136.5 50 139.5 ;
      LAYER METG1 ;
        RECT 0 136.5 50 139.5 ;
      LAYER METS2 ;
        RECT 0 136.5 50 139.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 152.5 50 155.5 ;
      LAYER METG1 ;
        RECT 0 152.5 50 155.5 ;
      LAYER METS2 ;
        RECT 0 152.5 50 155.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 156.5 50 159.5 ;
      LAYER METG1 ;
        RECT 0 156.5 50 159.5 ;
      LAYER METS2 ;
        RECT 0 156.5 50 159.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 160.5 50 163.5 ;
      LAYER METG1 ;
        RECT 0 160.5 50 163.5 ;
      LAYER METS2 ;
        RECT 0 160.5 50 163.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET6 ;
        RECT 0 4.5 50 7.5 ;
      LAYER METG1 ;
        RECT 0 4.5 50 7.5 ;
      LAYER METS2 ;
        RECT 0 4.5 50 7.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 8.5 50 11.5 ;
      LAYER METG1 ;
        RECT 0 8.5 50 11.5 ;
      LAYER METS2 ;
        RECT 0 8.5 50 11.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 20.5 50 23.5 ;
      LAYER METG1 ;
        RECT 0 20.5 50 23.5 ;
      LAYER METS2 ;
        RECT 0 20.5 50 23.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 24.5 50 27.5 ;
      LAYER METG1 ;
        RECT 0 24.5 50 27.5 ;
      LAYER METS2 ;
        RECT 0 24.5 50 27.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 36.5 50 39.5 ;
      LAYER METG1 ;
        RECT 0 36.5 50 39.5 ;
      LAYER METS2 ;
        RECT 0 36.5 50 39.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 44.5 50 47.5 ;
      LAYER METG1 ;
        RECT 0 44.5 50 47.5 ;
      LAYER METS2 ;
        RECT 0 44.5 50 47.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 52.5 50 55.5 ;
      LAYER METG1 ;
        RECT 0 52.5 50 55.5 ;
      LAYER METS2 ;
        RECT 0 52.5 50 55.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 60.5 50 63.5 ;
      LAYER METG1 ;
        RECT 0 60.5 50 63.5 ;
      LAYER METS2 ;
        RECT 0 60.5 50 63.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 68.5 50 71.5 ;
      LAYER METG1 ;
        RECT 0 68.5 50 71.5 ;
      LAYER METS2 ;
        RECT 0 68.5 50 71.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 100.5 50 103.5 ;
      LAYER METG1 ;
        RECT 0 100.5 50 103.5 ;
      LAYER METS2 ;
        RECT 0 100.5 50 103.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 104.5 50 107.5 ;
      LAYER METG1 ;
        RECT 0 104.5 50 107.5 ;
      LAYER METS2 ;
        RECT 0 104.5 50 107.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 112.5 50 115.5 ;
      LAYER METG1 ;
        RECT 0 112.5 50 115.5 ;
      LAYER METS2 ;
        RECT 0 112.5 50 115.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 116.5 50 119.5 ;
      LAYER METG1 ;
        RECT 0 116.5 50 119.5 ;
      LAYER METS2 ;
        RECT 0 116.5 50 119.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 120.5 50 123.5 ;
      LAYER METG1 ;
        RECT 0 120.5 50 123.5 ;
      LAYER METS2 ;
        RECT 0 120.5 50 123.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 124.5 50 127.5 ;
      LAYER METG1 ;
        RECT 0 124.5 50 127.5 ;
      LAYER METS2 ;
        RECT 0 124.5 50 127.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 132.5 50 135.5 ;
      LAYER METG1 ;
        RECT 0 132.5 50 135.5 ;
      LAYER METS2 ;
        RECT 0 132.5 50 135.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 140.5 50 143.5 ;
      LAYER METG1 ;
        RECT 0 140.5 50 143.5 ;
      LAYER METS2 ;
        RECT 0 140.5 50 143.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 144.5 50 147.5 ;
      LAYER METG1 ;
        RECT 0 144.5 50 147.5 ;
      LAYER METS2 ;
        RECT 0 144.5 50 147.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 148.5 50 151.5 ;
      LAYER METG1 ;
        RECT 0 148.5 50 151.5 ;
      LAYER METS2 ;
        RECT 0 148.5 50 151.5 ;
    END
  END VSS
  OBS
    LAYER CUT56 ;
      RECT 0 0 50 170 ;
    LAYER MET6 ;
      RECT 0 0 50 170 ;
    LAYER CUTS1 ;
      RECT 0 0 50 170 ;
    LAYER METS1 ;
      RECT 0 0 50 170 ;
    LAYER CUTS2 ;
      RECT 0 0 50 170 ;
    LAYER METS2 ;
      RECT 0 0 50 170 ;
    LAYER CUTS3 ;
      RECT 0 0 50 170 ;
    LAYER METS3 ;
      RECT 0 0 50 170 ;
    LAYER CUTG1 ;
      RECT 0 0 50 170 ;
    LAYER METG1 ;
      RECT 0 0 50 170 ;
    LAYER CUTG2 ;
      RECT 0 0 50 170 ;
    LAYER METG2 ;
      RECT 0 0 50 170 ;
    LAYER CUTTOP ;
      RECT 0 0 50 170 ;
    LAYER METTOP ;
      RECT 0 0 50 170 ;
      LAYER OVLAP ;
       RECT 0.000 84.000 50.000 86.000 ;
  END
END IOCB2EWDA5C0A1


MACRO IOCB2EWGA5C0A1
  CLASS PAD POWER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EWGA5C0A1 0 0 ;
  SIZE 50 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET6 ;
        RECT 0 12.5 50 15.5 ;
      LAYER METG1 ;
        RECT 0 12.5 50 15.5 ;
      LAYER METS2 ;
        RECT 0 12.5 50 15.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 16.5 50 19.5 ;
      LAYER METG1 ;
        RECT 0 16.5 50 19.5 ;
      LAYER METS2 ;
        RECT 0 16.5 50 19.5 ;
    END
  END VDD
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET6 ;
        RECT 0 28.5 50 31.5 ;
      LAYER METG1 ;
        RECT 0 28.5 50 31.5 ;
      LAYER METS2 ;
        RECT 0 28.5 50 31.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 32.5 50 35.5 ;
      LAYER METG1 ;
        RECT 0 32.5 50 35.5 ;
      LAYER METS2 ;
        RECT 0 32.5 50 35.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 40.5 50 43.5 ;
      LAYER METG1 ;
        RECT 0 40.5 50 43.5 ;
      LAYER METS2 ;
        RECT 0 40.5 50 43.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 48.5 50 51.5 ;
      LAYER METG1 ;
        RECT 0 48.5 50 51.5 ;
      LAYER METS2 ;
        RECT 0 48.5 50 51.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 56.5 50 59.5 ;
      LAYER METG1 ;
        RECT 0 56.5 50 59.5 ;
      LAYER METS2 ;
        RECT 0 56.5 50 59.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 64.5 50 67.5 ;
      LAYER METG1 ;
        RECT 0 64.5 50 67.5 ;
      LAYER METS2 ;
        RECT 0 64.5 50 67.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 72.5 50 75.5 ;
      LAYER METG1 ;
        RECT 0 72.5 50 75.5 ;
      LAYER METS2 ;
        RECT 0 72.5 50 75.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 76.5 50 79.5 ;
      LAYER METG1 ;
        RECT 0 76.5 50 79.5 ;
      LAYER METS2 ;
        RECT 0 76.5 50 79.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 80.5 50 83.5 ;
      LAYER METG1 ;
        RECT 0 80.5 50 83.5 ;
      LAYER METS2 ;
        RECT 0 80.5 50 83.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 84.5 50 87.5 ;
      LAYER METG1 ;
        RECT 0 84.5 50 87.5 ;
      LAYER METS2 ;
        RECT 0 84.5 50 87.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 88.5 50 91.5 ;
      LAYER METG1 ;
        RECT 0 88.5 50 91.5 ;
      LAYER METS2 ;
        RECT 0 88.5 50 91.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 92.5 50 95.5 ;
      LAYER METG1 ;
        RECT 0 92.5 50 95.5 ;
      LAYER METS2 ;
        RECT 0 92.5 50 95.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 96.5 50 99.5 ;
      LAYER METG1 ;
        RECT 0 96.5 50 99.5 ;
      LAYER METS2 ;
        RECT 0 96.5 50 99.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 108.5 50 111.5 ;
      LAYER METG1 ;
        RECT 0 108.5 50 111.5 ;
      LAYER METS2 ;
        RECT 0 108.5 50 111.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 128.5 50 131.5 ;
      LAYER METG1 ;
        RECT 0 128.5 50 131.5 ;
      LAYER METS2 ;
        RECT 0 128.5 50 131.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 136.5 50 139.5 ;
      LAYER METG1 ;
        RECT 0 136.5 50 139.5 ;
      LAYER METS2 ;
        RECT 0 136.5 50 139.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 152.5 50 155.5 ;
      LAYER METG1 ;
        RECT 0 152.5 50 155.5 ;
      LAYER METS2 ;
        RECT 0 152.5 50 155.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 156.5 50 159.5 ;
      LAYER METG1 ;
        RECT 0 156.5 50 159.5 ;
      LAYER METS2 ;
        RECT 0 156.5 50 159.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 160.5 50 163.5 ;
      LAYER METG1 ;
        RECT 0 160.5 50 163.5 ;
      LAYER METS2 ;
        RECT 0 160.5 50 163.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET6 ;
        RECT 0 4.5 50 7.5 ;
      LAYER METG1 ;
        RECT 0 4.5 50 7.5 ;
      LAYER METS2 ;
        RECT 0 4.5 50 7.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 8.5 50 11.5 ;
      LAYER METG1 ;
        RECT 0 8.5 50 11.5 ;
      LAYER METS2 ;
        RECT 0 8.5 50 11.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 20.5 50 23.5 ;
      LAYER METG1 ;
        RECT 0 20.5 50 23.5 ;
      LAYER METS2 ;
        RECT 0 20.5 50 23.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 24.5 50 27.5 ;
      LAYER METG1 ;
        RECT 0 24.5 50 27.5 ;
      LAYER METS2 ;
        RECT 0 24.5 50 27.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 36.5 50 39.5 ;
      LAYER METG1 ;
        RECT 0 36.5 50 39.5 ;
      LAYER METS2 ;
        RECT 0 36.5 50 39.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 44.5 50 47.5 ;
      LAYER METG1 ;
        RECT 0 44.5 50 47.5 ;
      LAYER METS2 ;
        RECT 0 44.5 50 47.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 52.5 50 55.5 ;
      LAYER METG1 ;
        RECT 0 52.5 50 55.5 ;
      LAYER METS2 ;
        RECT 0 52.5 50 55.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 60.5 50 63.5 ;
      LAYER METG1 ;
        RECT 0 60.5 50 63.5 ;
      LAYER METS2 ;
        RECT 0 60.5 50 63.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 68.5 50 71.5 ;
      LAYER METG1 ;
        RECT 0 68.5 50 71.5 ;
      LAYER METS2 ;
        RECT 0 68.5 50 71.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 100.5 50 103.5 ;
      LAYER METG1 ;
        RECT 0 100.5 50 103.5 ;
      LAYER METS2 ;
        RECT 0 100.5 50 103.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 104.5 50 107.5 ;
      LAYER METG1 ;
        RECT 0 104.5 50 107.5 ;
      LAYER METS2 ;
        RECT 0 104.5 50 107.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 112.5 50 115.5 ;
      LAYER METG1 ;
        RECT 0 112.5 50 115.5 ;
      LAYER METS2 ;
        RECT 0 112.5 50 115.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 116.5 50 119.5 ;
      LAYER METG1 ;
        RECT 0 116.5 50 119.5 ;
      LAYER METS2 ;
        RECT 0 116.5 50 119.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 120.5 50 123.5 ;
      LAYER METG1 ;
        RECT 0 120.5 50 123.5 ;
      LAYER METS2 ;
        RECT 0 120.5 50 123.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 124.5 50 127.5 ;
      LAYER METG1 ;
        RECT 0 124.5 50 127.5 ;
      LAYER METS2 ;
        RECT 0 124.5 50 127.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 132.5 50 135.5 ;
      LAYER METG1 ;
        RECT 0 132.5 50 135.5 ;
      LAYER METS2 ;
        RECT 0 132.5 50 135.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 140.5 50 143.5 ;
      LAYER METG1 ;
        RECT 0 140.5 50 143.5 ;
      LAYER METS2 ;
        RECT 0 140.5 50 143.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 144.5 50 147.5 ;
      LAYER METG1 ;
        RECT 0 144.5 50 147.5 ;
      LAYER METS2 ;
        RECT 0 144.5 50 147.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 148.5 50 151.5 ;
      LAYER METG1 ;
        RECT 0 148.5 50 151.5 ;
      LAYER METS2 ;
        RECT 0 148.5 50 151.5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG2 ;
        RECT 14.5 0 20.5 5 ;
      LAYER METTOP ;
        RECT 14.5 0 20.5 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG2 ;
        RECT 22 0 28 5 ;
      LAYER METTOP ;
        RECT 22 0 28 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG2 ;
        RECT 29.5 0 35.5 5 ;
      LAYER METTOP ;
        RECT 29.5 0 35.5 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG2 ;
        RECT 37 0 43 5 ;
      LAYER METTOP ;
        RECT 37 0 43 5 ;
    END
    PORT
      CLASS CORE ;
      LAYER METG2 ;
        RECT 7 0 13 5 ;
      LAYER METTOP ;
        RECT 7 0 13 5 ;
    END
  END VSS
  OBS
    LAYER CUT56 ;
      RECT 0 0 50 170 ;
    LAYER MET6 ;
      RECT 0 0 50 170 ;
    LAYER CUTS1 ;
      RECT 0 0 50 170 ;
    LAYER METS1 ;
      RECT 0 0 50 170 ;
    LAYER CUTS2 ;
      RECT 0 0 50 170 ;
    LAYER METS2 ;
      RECT 0 0 50 170 ;
    LAYER CUTS3 ;
      RECT 0 0 50 170 ;
    LAYER METS3 ;
      RECT 0 0 50 170 ;
    LAYER CUTG1 ;
      RECT 0 0 50 170 ;
    LAYER METG1 ;
      RECT 0 0 50 170 ;
    LAYER CUTG2 ;
      RECT 0 0 50 170 ;
    LAYER METG2 ;
      RECT 0 0 50 170 ;
    LAYER CUTTOP ;
      RECT 0 0 50 170 ;
    LAYER METTOP ;
      RECT 0 0 50 170 ;
      LAYER OVLAP ;
       RECT 0.000 84.000 50.000 86.000 ;
  END
END IOCB2EWGA5C0A1


MACRO IOCB2EWSA5C0A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN IOCB2EWSA5C0A1 0 0 ;
  SIZE 40 BY 170 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE170 ;
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET6 ;
        RECT 0 12.5 40 15.5 ;
      LAYER METG1 ;
        RECT 0 12.5 40 15.5 ;
      LAYER METS1 ;
        RECT 0 12.5 40 15.5 ;
      LAYER METS2 ;
        RECT 0 12.5 40 15.5 ;
      LAYER METS3 ;
        RECT 0 12.5 40 15.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 16.5 40 19.5 ;
      LAYER METG1 ;
        RECT 0 16.5 40 19.5 ;
      LAYER METS1 ;
        RECT 0 16.5 40 19.5 ;
      LAYER METS2 ;
        RECT 0 16.5 40 19.5 ;
      LAYER METS3 ;
        RECT 0 16.5 40 19.5 ;
    END
  END VDD
  PIN VDE
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET6 ;
        RECT 0 28.5 40 31.5 ;
      LAYER METG1 ;
        RECT 0 28.5 40 31.5 ;
      LAYER METS1 ;
        RECT 0 28.5 40 31.5 ;
      LAYER METS2 ;
        RECT 0 28.5 40 31.5 ;
      LAYER METS3 ;
        RECT 0 28.5 40 31.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 32.5 40 35.5 ;
      LAYER METG1 ;
        RECT 0 32.5 40 35.5 ;
      LAYER METS1 ;
        RECT 0 32.5 40 35.5 ;
      LAYER METS2 ;
        RECT 0 32.5 40 35.5 ;
      LAYER METS3 ;
        RECT 0 32.5 40 35.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 40.5 40 43.5 ;
      LAYER METG1 ;
        RECT 0 40.5 40 43.5 ;
      LAYER METS1 ;
        RECT 0 40.5 40 43.5 ;
      LAYER METS2 ;
        RECT 0 40.5 40 43.5 ;
      LAYER METS3 ;
        RECT 0 40.5 40 43.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 48.5 40 51.5 ;
      LAYER METG1 ;
        RECT 0 48.5 40 51.5 ;
      LAYER METS1 ;
        RECT 0 48.5 40 51.5 ;
      LAYER METS2 ;
        RECT 0 48.5 40 51.5 ;
      LAYER METS3 ;
        RECT 0 48.5 40 51.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 56.5 40 59.5 ;
      LAYER METG1 ;
        RECT 0 56.5 40 59.5 ;
      LAYER METS1 ;
        RECT 0 56.5 40 59.5 ;
      LAYER METS2 ;
        RECT 0 56.5 40 59.5 ;
      LAYER METS3 ;
        RECT 0 56.5 40 59.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 64.5 40 67.5 ;
      LAYER METG1 ;
        RECT 0 64.5 40 67.5 ;
      LAYER METS1 ;
        RECT 0 64.5 40 67.5 ;
      LAYER METS2 ;
        RECT 0 64.5 40 67.5 ;
      LAYER METS3 ;
        RECT 0 64.5 40 67.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 72.5 40 75.5 ;
      LAYER METG1 ;
        RECT 0 72.5 40 75.5 ;
      LAYER METS1 ;
        RECT 0 72.5 40 75.5 ;
      LAYER METS2 ;
        RECT 0 72.5 40 75.5 ;
      LAYER METS3 ;
        RECT 0 72.5 40 75.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 76.5 40 79.5 ;
      LAYER METG1 ;
        RECT 0 76.5 40 79.5 ;
      LAYER METS1 ;
        RECT 0 76.5 40 79.5 ;
      LAYER METS2 ;
        RECT 0 76.5 40 79.5 ;
      LAYER METS3 ;
        RECT 0 76.5 40 79.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 80.5 40 83.5 ;
      LAYER METG1 ;
        RECT 0 80.5 40 83.5 ;
      LAYER METS1 ;
        RECT 0 80.5 40 83.5 ;
      LAYER METS2 ;
        RECT 0 80.5 40 83.5 ;
      LAYER METS3 ;
        RECT 0 80.5 40 83.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 84.5 40 87.5 ;
      LAYER METG1 ;
        RECT 0 84.5 40 87.5 ;
      LAYER METS1 ;
        RECT 0 84.5 40 87.5 ;
      LAYER METS2 ;
        RECT 0 84.5 40 87.5 ;
      LAYER METS3 ;
        RECT 0 84.5 40 87.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 88.5 40 91.5 ;
      LAYER METG1 ;
        RECT 0 88.5 40 91.5 ;
      LAYER METS1 ;
        RECT 0 88.5 40 91.5 ;
      LAYER METS2 ;
        RECT 0 88.5 40 91.5 ;
      LAYER METS3 ;
        RECT 0 88.5 40 91.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 92.5 40 95.5 ;
      LAYER METG1 ;
        RECT 0 92.5 40 95.5 ;
      LAYER METS1 ;
        RECT 0 92.5 40 95.5 ;
      LAYER METS2 ;
        RECT 0 92.5 40 95.5 ;
      LAYER METS3 ;
        RECT 0 92.5 40 95.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 96.5 40 99.5 ;
      LAYER METG1 ;
        RECT 0 96.5 40 99.5 ;
      LAYER METS1 ;
        RECT 0 96.5 40 99.5 ;
      LAYER METS2 ;
        RECT 0 96.5 40 99.5 ;
      LAYER METS3 ;
        RECT 0 96.5 40 99.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 108.5 40 111.5 ;
      LAYER METG1 ;
        RECT 0 108.5 40 111.5 ;
      LAYER METS1 ;
        RECT 0 108.5 40 111.5 ;
      LAYER METS2 ;
        RECT 0 108.5 40 111.5 ;
      LAYER METS3 ;
        RECT 0 108.5 40 111.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 128.5 40 131.5 ;
      LAYER METG1 ;
        RECT 0 128.5 40 131.5 ;
      LAYER METS1 ;
        RECT 0 128.5 40 131.5 ;
      LAYER METS2 ;
        RECT 0 128.5 40 131.5 ;
      LAYER METS3 ;
        RECT 0 128.5 40 131.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 136.5 40 139.5 ;
      LAYER METG1 ;
        RECT 0 136.5 40 139.5 ;
      LAYER METS1 ;
        RECT 0 136.5 40 139.5 ;
      LAYER METS2 ;
        RECT 0 136.5 40 139.5 ;
      LAYER METS3 ;
        RECT 0 136.5 40 139.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 152.5 40 155.5 ;
      LAYER METG1 ;
        RECT 0 152.5 40 155.5 ;
      LAYER METS1 ;
        RECT 0 152.5 40 155.5 ;
      LAYER METS2 ;
        RECT 0 152.5 40 155.5 ;
      LAYER METS3 ;
        RECT 0 152.5 40 155.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 156.5 40 159.5 ;
      LAYER METG1 ;
        RECT 0 156.5 40 159.5 ;
      LAYER METS1 ;
        RECT 0 156.5 40 159.5 ;
      LAYER METS2 ;
        RECT 0 156.5 40 159.5 ;
      LAYER METS3 ;
        RECT 0 156.5 40 159.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 160.5 40 163.5 ;
      LAYER METG1 ;
        RECT 0 160.5 40 163.5 ;
      LAYER METS1 ;
        RECT 0 160.5 40 163.5 ;
      LAYER METS2 ;
        RECT 0 160.5 40 163.5 ;
      LAYER METS3 ;
        RECT 0 160.5 40 163.5 ;
    END
  END VDE
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE FEEDTHRU ;
    PORT
      LAYER MET6 ;
        RECT 0 4.5 40 7.5 ;
      LAYER METG1 ;
        RECT 0 4.5 40 7.5 ;
      LAYER METS1 ;
        RECT 0 4.5 40 7.5 ;
      LAYER METS2 ;
        RECT 0 4.5 40 7.5 ;
      LAYER METS3 ;
        RECT 0 4.5 40 7.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 8.5 40 11.5 ;
      LAYER METG1 ;
        RECT 0 8.5 40 11.5 ;
      LAYER METS1 ;
        RECT 0 8.5 40 11.5 ;
      LAYER METS2 ;
        RECT 0 8.5 40 11.5 ;
      LAYER METS3 ;
        RECT 0 8.5 40 11.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 20.5 40 23.5 ;
      LAYER METG1 ;
        RECT 0 20.5 40 23.5 ;
      LAYER METS1 ;
        RECT 0 20.5 40 23.5 ;
      LAYER METS2 ;
        RECT 0 20.5 40 23.5 ;
      LAYER METS3 ;
        RECT 0 20.5 40 23.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 24.5 40 27.5 ;
      LAYER METG1 ;
        RECT 0 24.5 40 27.5 ;
      LAYER METS1 ;
        RECT 0 24.5 40 27.5 ;
      LAYER METS2 ;
        RECT 0 24.5 40 27.5 ;
      LAYER METS3 ;
        RECT 0 24.5 40 27.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 36.5 40 39.5 ;
      LAYER METG1 ;
        RECT 0 36.5 40 39.5 ;
      LAYER METS1 ;
        RECT 0 36.5 40 39.5 ;
      LAYER METS2 ;
        RECT 0 36.5 40 39.5 ;
      LAYER METS3 ;
        RECT 0 36.5 40 39.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 44.5 40 47.5 ;
      LAYER METG1 ;
        RECT 0 44.5 40 47.5 ;
      LAYER METS1 ;
        RECT 0 44.5 40 47.5 ;
      LAYER METS2 ;
        RECT 0 44.5 40 47.5 ;
      LAYER METS3 ;
        RECT 0 44.5 40 47.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 52.5 40 55.5 ;
      LAYER METG1 ;
        RECT 0 52.5 40 55.5 ;
      LAYER METS1 ;
        RECT 0 52.5 40 55.5 ;
      LAYER METS2 ;
        RECT 0 52.5 40 55.5 ;
      LAYER METS3 ;
        RECT 0 52.5 40 55.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 60.5 40 63.5 ;
      LAYER METG1 ;
        RECT 0 60.5 40 63.5 ;
      LAYER METS1 ;
        RECT 0 60.5 40 63.5 ;
      LAYER METS2 ;
        RECT 0 60.5 40 63.5 ;
      LAYER METS3 ;
        RECT 0 60.5 40 63.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 68.5 40 71.5 ;
      LAYER METG1 ;
        RECT 0 68.5 40 71.5 ;
      LAYER METS1 ;
        RECT 0 68.5 40 71.5 ;
      LAYER METS2 ;
        RECT 0 68.5 40 71.5 ;
      LAYER METS3 ;
        RECT 0 68.5 40 71.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 100.5 40 103.5 ;
      LAYER METG1 ;
        RECT 0 100.5 40 103.5 ;
      LAYER METS1 ;
        RECT 0 100.5 40 103.5 ;
      LAYER METS2 ;
        RECT 0 100.5 40 103.5 ;
      LAYER METS3 ;
        RECT 0 100.5 40 103.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 104.5 40 107.5 ;
      LAYER METG1 ;
        RECT 0 104.5 40 107.5 ;
      LAYER METS1 ;
        RECT 0 104.5 40 107.5 ;
      LAYER METS2 ;
        RECT 0 104.5 40 107.5 ;
      LAYER METS3 ;
        RECT 0 104.5 40 107.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 112.5 40 115.5 ;
      LAYER METG1 ;
        RECT 0 112.5 40 115.5 ;
      LAYER METS1 ;
        RECT 0 112.5 40 115.5 ;
      LAYER METS2 ;
        RECT 0 112.5 40 115.5 ;
      LAYER METS3 ;
        RECT 0 112.5 40 115.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 116.5 40 119.5 ;
      LAYER METG1 ;
        RECT 0 116.5 40 119.5 ;
      LAYER METS1 ;
        RECT 0 116.5 40 119.5 ;
      LAYER METS2 ;
        RECT 0 116.5 40 119.5 ;
      LAYER METS3 ;
        RECT 0 116.5 40 119.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 120.5 40 123.5 ;
      LAYER METG1 ;
        RECT 0 120.5 40 123.5 ;
      LAYER METS1 ;
        RECT 0 120.5 40 123.5 ;
      LAYER METS2 ;
        RECT 0 120.5 40 123.5 ;
      LAYER METS3 ;
        RECT 0 120.5 40 123.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 124.5 40 127.5 ;
      LAYER METG1 ;
        RECT 0 124.5 40 127.5 ;
      LAYER METS1 ;
        RECT 0 124.5 40 127.5 ;
      LAYER METS2 ;
        RECT 0 124.5 40 127.5 ;
      LAYER METS3 ;
        RECT 0 124.5 40 127.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 132.5 40 135.5 ;
      LAYER METG1 ;
        RECT 0 132.5 40 135.5 ;
      LAYER METS1 ;
        RECT 0 132.5 40 135.5 ;
      LAYER METS2 ;
        RECT 0 132.5 40 135.5 ;
      LAYER METS3 ;
        RECT 0 132.5 40 135.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 140.5 40 143.5 ;
      LAYER METG1 ;
        RECT 0 140.5 40 143.5 ;
      LAYER METS1 ;
        RECT 0 140.5 40 143.5 ;
      LAYER METS2 ;
        RECT 0 140.5 40 143.5 ;
      LAYER METS3 ;
        RECT 0 140.5 40 143.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 144.5 40 147.5 ;
      LAYER METG1 ;
        RECT 0 144.5 40 147.5 ;
      LAYER METS1 ;
        RECT 0 144.5 40 147.5 ;
      LAYER METS2 ;
        RECT 0 144.5 40 147.5 ;
      LAYER METS3 ;
        RECT 0 144.5 40 147.5 ;
    END
    PORT
      LAYER MET6 ;
        RECT 0 148.5 40 151.5 ;
      LAYER METG1 ;
        RECT 0 148.5 40 151.5 ;
      LAYER METS1 ;
        RECT 0 148.5 40 151.5 ;
      LAYER METS2 ;
        RECT 0 148.5 40 151.5 ;
      LAYER METS3 ;
        RECT 0 148.5 40 151.5 ;
    END
  END VSS
  OBS
    LAYER CUT56 ;
      RECT 0 0 40 170 ;
    LAYER MET6 ;
      RECT 0 0 40 170 ;
    LAYER CUTS1 ;
      RECT 0 0 40 170 ;
    LAYER METS1 ;
      RECT 0 0 40 170 ;
    LAYER CUTS2 ;
      RECT 0 0 40 170 ;
    LAYER METS2 ;
      RECT 0 0 40 170 ;
    LAYER CUTS3 ;
      RECT 0 0 40 170 ;
    LAYER METS3 ;
      RECT 0 0 40 170 ;
    LAYER CUTG1 ;
      RECT 0 0 40 170 ;
    LAYER METG1 ;
      RECT 0 0 40 170 ;
    LAYER CUTG2 ;
      RECT 0 0 40 170 ;
    LAYER METG2 ;
      RECT 0 0 40 170 ;
    LAYER CUTTOP ;
      RECT 0 0 40 170 ;
    LAYER METTOP ;
      RECT 0 0 40 170 ;
      LAYER OVLAP ;
       RECT 0.000 84.000 40.000 86.000 ;
  END
END IOCB2EWSA5C0A1


MACRO EXTGFCB2E25XC0A0
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN EXTGFCB2E25XC0A0 0 0 ;
  SIZE 48 BY 141 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE141 ;
  OBS
    LAYER METG2 ;
      RECT 0 0 48 141 ;
    LAYER CUTTOP ;
      RECT 0 0 48 141 ;
    LAYER METTOP ;
      RECT 0 0 48 141 ;
      LAYER OVLAP ;
       RECT 0.000 139.000 48.000 141.000 ;
  END
END EXTGFCB2E25XC0A0


#----------------------------------------------------------------
# Comment  : PAD Cell for 60um 
#----------------------------------------------------------------

MACRO EXTGOCB0316X70A1
  CLASS PAD SPACER ;
  ORIGIN 0 0 ;
  FOREIGN EXTGOCB0316X70A1 0 0 ;
  SIZE 40 BY 10 ;
  SYMMETRY X Y R90 ;
  SITE IOSITE10 ;
  OBS
    LAYER MET1 ;
      RECT -9 10 49 137 ;
    LAYER CUT12 ;
      RECT -9 10 49 137 ;
    LAYER MET2 ;
      RECT -9 10 49 137 ;
    LAYER CUT23 ;
      RECT -9 10 49 137 ;
    LAYER MET3 ;
      RECT -9 10 49 137 ;
    LAYER CUT34 ;
      RECT -9 10 49 137 ;
    LAYER MET4 ;
      RECT -9 10 49 137 ;
    LAYER CUT45 ;
      RECT -9 10 49 137 ;
    LAYER MET5 ;
      RECT -9 10 49 137 ;
    LAYER CUT56 ;
      RECT -9 10 49 137 ;
    LAYER MET6 ;
      RECT -9 10 49 137 ;
    LAYER CUTS1 ;
      RECT -9 10 49 137 ;
    LAYER METS1 ;
      RECT -9 10 49 137 ;
    LAYER CUTS2 ;
      RECT -9 10 49 137 ;
    LAYER METS2 ;
      RECT -9 10 49 137 ;
    LAYER CUTS3 ;
      RECT -9 10 49 137 ;
    LAYER METS3 ;
      RECT -9 10 49 137 ;
    LAYER CUTS4 ;
      RECT -9 10 49 137 ;
    LAYER METS4 ;
      RECT -9 10 49 137 ;
    LAYER CUTG1 ;
      RECT -9 10 49 137 ;
    LAYER METG1 ;
      RECT -9 10 49 137 ;
    LAYER CUTG2 ;
      RECT -9 10 49 137 ;
    LAYER METG2 ;
      RECT -9 10 49 137 ;
    LAYER CUTTOP ;
      RECT -9 10 49 137 ;
    LAYER METTOP ;
      RECT -9 10 49 137 ;
      LAYER OVLAP ;
       RECT 0.000 8.000 40.000 10.000 ;
  END
END EXTGOCB0316X70A1


#----- CS202 Monitor LEF ---------------------------------------------
# Rev0001 07/06/15 : New Release(FrameSize=100x100um)          C.Sato
#                     (for 50I_STD)
#---------------------------------------------------------------------
#--- CS202 CORNER MONITOR CELL LEF ----------------------------------
#----- 50umInline(50I_STD) ---------------------------
MACRO ZMGACS202S_50I
  CLASS ENDCAP TOPRIGHT ;
  ORIGIN 0 0 ;
  FOREIGN ZMGACS202S_50I 0 0 ;
  SIZE 100 BY 100 ;
  SYMMETRY X Y R90 ;
   OBS
      LAYER OVLAP ;
       RECT 98.000 98.000 100.000 100.000 ;
   END
END ZMGACS202S_50I


MACRO ZMGBCS202S_50I
  CLASS ENDCAP TOPLEFT ;
  ORIGIN 0 0 ;
  FOREIGN ZMGBCS202S_50I 0 0 ;
  SIZE 100 BY 100 ;
  SYMMETRY X Y R90 ;
   OBS
      LAYER OVLAP ;
       RECT 98.000 98.000 100.000 100.000 ;
   END
END ZMGBCS202S_50I


MACRO ZMGCCS202S_50I
  CLASS ENDCAP BOTTOMLEFT ;
  ORIGIN 0 0 ;
  FOREIGN ZMGCCS202S_50I 0 0 ;
  SIZE 100 BY 100 ;
  SYMMETRY X Y R90 ;
   OBS
      LAYER OVLAP ;
       RECT 98.000 98.000 100.000 100.000 ;
   END
END ZMGCCS202S_50I


MACRO ZMGDCS202S_50I
  CLASS ENDCAP BOTTOMRIGHT ;
  ORIGIN 0 0 ;
  FOREIGN ZMGDCS202S_50I 0 0 ;
  SIZE 100 BY 100 ;
  SYMMETRY X Y R90 ;
   OBS
      LAYER OVLAP ;
       RECT 98.000 98.000 100.000 100.000 ;
   END
END ZMGDCS202S_50I
#--------------------------------------------------------------------
END LIBRARY
# FUJITSU MICROELECTRONICS Proprietary and Confidential
#-----------------------------------------------------------------------
# Technology rule (65nm S/C LEF FOR 7LAYER ROUTING - LEF5.6)
#                       CS200L PROCESS
#-----------------------------------------------------------------------
#
#  [Layers Information of 7layer]
#     #layer    layerName   pitch   width   spacing   direction
#     layer7     METTOP     1.60    0.80    0.80      H
#     layer6     METG1      0.80    0.40    0.40      V
#     layer5     MET5       0.20    0.10    0.10      H
#     layer4     MET4       0.20    0.10    0.10      V
#     layer3     MET3       0.20    0.10    0.10      H
#     layer2     MET2       0.20    0.10    0.10      V
#     layer1     MET1       0.20    0.10    0.10      H
#
#  [Structure] RF_METAL : 7S0G1
#     metal1
#     intermediate metal1 - intermediate metal4
#     global metal1
#     top metal
#
#  [History]
#   o Revision 004 07/02/2008
#      Reference document
#       - CS200L DESIGN RULE REVISION 2.1
#      Additional Rule
#       - The spacing rule more than the width of 100um is changed.(0.80um->1.12um)
#   o Revision 003 04/02/2008
#      Reference document
#       - CS200L DESIGN RULE REVISION 1.2
#       - CS200A DESIGN RULE REVISION 1.8
#      Additional Rule
#       - VIA-Fig(Double VIA/Triple VIA/Asymmetric single VIA) are added
#       - PWELL/NWELL Layer are added
#   o Revision 002 05/31/2007
#      Reference document
#       - CS200L DESIGN RULE REVISION 1.0
#       - CS200A DESIGN RULE REVISION 1.62
#      Additional Rule
#       - NONDEFAULTRULE(WIDEWIRE/WIDEWIRE_DC) are added
#       - VIA-Fig(VIA34P2/VIA1_2NV/VIA1_2SV) are added
#   o Revision 001 06/26/2006
#      Reference document
#       - CS200A DESIGN RULE REVISION 1.3
#
#  [Release Note]
#   o Resistance and capacity must use the capacity table prepared with each tool.
#         First Encounter : Capacitance Table File
#         PhyC, Astro     : TLU+
#   o Spacing rule for high voltage(1.8v/2.5v/3.3v) cannot be treated on LEF.
#     Please do not use the wiring for high voltage(1.8v/2.5v/3.3v) in the core area.
#   o The wiring for 45 degrees is not supported.
#
#  [Designer]
#     M.Sekido
#
#-----------------------------------------------------------------------
# Copyright (c) 2006-2008 FUJITSU MICROELECTRONICS LIMITED All rights reserved.
#

VERSION 5.6 ;
# === LEF v5.5 SPEC ===
#NAMESCASESENSITIVE ON ;
# === END ===
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;
USEMINSPACING OBS OFF ;
# === LEF v5.5 SPEC ===
#USEMINSPACING PIN OFF ;
# === END ===
CLEARANCEMEASURE EUCLIDEAN ;

# === LEF v5.6 SPEC ===
PROPERTYDEFINITIONS
  LAYER LEF57_ENCLOSURE STRING ;
  LAYER LEF57_MINSTEP STRING ;
  LAYER LEF57_ANTENNACUMROUTINGPLUSCUT STRING ;
  LAYER LEF57_ANTENNAAREAMINUSDIFF STRING ;
  LAYER LEF58_TYPE STRING ;
  LAYER LEF57_SPACING STRING ;
  LAYER LEF58_WIDTH STRING ;
  LAYER LEF58_VOLTAGESPACING STRING ;
END PROPERTYDEFINITIONS
# === END ===

#  ANTENNAINPUTGATEAREA  0.0840 ;
#  ANTENNAINOUTDIFFAREA  0.0231 ;
#  ANTENNAOUTPUTDIFFAREA 0.0231 ;

LAYER NWELL
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
  PROPERTY LEF58_WIDTH "WIDTH 0.44 ;" ;
#  PROPERTY LEF57_SPACING "SPACING 0.44 ;" ;
END NWELL

LAYER PWELL
  TYPE MASTERSLICE ;
  PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
#  PROPERTY LEF57_WIDTH "WIDTH 0.44 ;" ;
END PWELL

LAYER POLY
  TYPE MASTERSLICE ;
END POLY

LAYER DIFF
  TYPE MASTERSLICE ;
END DIFF

LAYER DIFFN
  TYPE MASTERSLICE ;
END DIFFN

LAYER DIFFP
  TYPE MASTERSLICE ;
END DIFFP

LAYER BUMPINH
  TYPE MASTERSLICE ;
END BUMPINH

LAYER BUMPIFS
  TYPE MASTERSLICE ;
END BUMPIFS

LAYER CUT78
  TYPE MASTERSLICE ;
END CUT78

LAYER MET8
  TYPE MASTERSLICE ;
END MET8

LAYER CUT67
  TYPE MASTERSLICE ;
END CUT67

LAYER MET7
  TYPE MASTERSLICE ;
END MET7

LAYER CUT56
  TYPE MASTERSLICE ;
END CUT56

LAYER MET6
  TYPE MASTERSLICE ;
END MET6

LAYER CUTS4
  TYPE MASTERSLICE ;
END CUTS4

LAYER METS4
  TYPE MASTERSLICE ;
END METS4

LAYER CUTS3
  TYPE MASTERSLICE ;
END CUTS3

LAYER METS3
  TYPE MASTERSLICE ;
END METS3

LAYER CUTS2
  TYPE MASTERSLICE ;
END CUTS2

LAYER METS2
  TYPE MASTERSLICE ;
END METS2

LAYER CUTS1
  TYPE MASTERSLICE ;
END CUTS1

LAYER METS1
  TYPE MASTERSLICE ;
END METS1

LAYER CUTG2
  TYPE MASTERSLICE ;
END CUTG2

LAYER METG2
  TYPE MASTERSLICE ;
END METG2

LAYER CUTT1
  TYPE MASTERSLICE ;
END CUTT1

LAYER METT1
  TYPE MASTERSLICE ;
END METT1

LAYER CUT01
  TYPE CUT ;
  SPACING 0.110 ;
END CUT01

LAYER MET1
  TYPE ROUTING ;
  PITCH 0.200 ;
  OFFSET 0.200 ;
  WIDTH 0.100 ;
  MINWIDTH 0.090 ;
  MAXWIDTH 3.000 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_MINSTEP "MINSTEP 0.045 MAXEDGES 1 ;" ;
# === END ===
  AREA 0.038 ;
  PROPERTY LEF58_VOLTAGESPACING "VOLTAGESPACING 0.9 0.1 5.0 0.3 ; VOLTAGESPACING TOCUT BELOW 0.9 0.1 5.0 0.5 ; VOLTAGESPACING TOCUT ABOVE 0.9 0.1 5.0 0.5 ;" ;
  MINENCLOSEDAREA 0.110 ;
  MINENCLOSEDAREA 0.800 WIDTH 0.210 ;
  MINENCLOSEDAREA 3.200 WIDTH 1.500 ;
  MINIMUMCUT 2 WIDTH 0.299 ;
  MINIMUMCUT 3 WIDTH 0.699 ;
  MINIMUMCUT 2 WIDTH 0.299 LENGTH 0.774 WITHIN 20000 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.000  0.180  0.380
    WIDTH 0.000        0.090  0.090  0.090
    WIDTH 0.150        0.100  0.120  0.120
    WIDTH 0.180        0.120  0.120  0.120
    WIDTH 0.210        0.120  0.120  0.150
    WIDTH 0.320        0.140  0.140  0.150
    WIDTH 1.500        0.140  0.140  0.500 ;
  MINIMUMDENSITY 20.000 ;
  MAXIMUMDENSITY 80.000 ;
  DENSITYCHECKWINDOW 40.000 40.000 ;
  DENSITYCHECKSTEP 10.000 ;
  DIRECTION HORIZONTAL ;
# === LEF v5.5 SPEC ===
#  ANTENNACUMAREARATIO 400.0 ;
#  ANTENNACUMDIFFAREARATIO PWL
#   ( ( 0.00000  400.0 ) ( 0.01919 400.0 ) ( 0.01920 100000.000 )
#     ( 1000.00000 100000.000 ) ) ;
#  ANTENNAAREAFACTOR 1.1 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_ANTENNACUMROUTINGPLUSCUT "ANTENNACUMROUTINGPLUSCUT ;" ;
  PROPERTY LEF57_ANTENNAAREAMINUSDIFF "ANTENNAAREAMINUSDIFF 118750 ;" ;
  ANTENNACUMDIFFAREARATIO 2000.0 ;
  ANTENNAAREAFACTOR 1.0 ;
# === END ===
END MET1

LAYER CUT12
  TYPE CUT ;
  SPACING 0.100 ;
# === LEF v5.6 SPEC ===
  ENCLOSURE BELOW 0.000 0.040 ;
  ENCLOSURE BELOW 0.015 0.040 WIDTH 0.501 ;
  ENCLOSURE BELOW 0.035 0.040 WIDTH 1.201 ;
  ENCLOSURE ABOVE 0.000 0.040 ;
  ENCLOSURE ABOVE 0.015 0.040 WIDTH 0.801 ;
  ENCLOSURE ABOVE 0.035 0.040 WIDTH 1.201 ;
# === END ===
# === LEF v5.5 SPEC ===
#  ANTENNACUMAREARATIO 1600.0 ;
#  ANTENNACUMDIFFAREARATIO PWL
#   ( ( 0.00000  1600.0 ) ( 0.01919 1600.0 ) ( 0.01920 100000.000 )
#     ( 1000.00000 100000.000 ) ) ;
#  ANTENNAAREAFACTOR 100.0 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_ANTENNACUMROUTINGPLUSCUT "ANTENNACUMROUTINGPLUSCUT ;" ;
  PROPERTY LEF57_ANTENNAAREAMINUSDIFF "ANTENNAAREAMINUSDIFF 118750 ;" ;
  ANTENNACUMDIFFAREARATIO 2000.0 ;
  ANTENNAAREAFACTOR 100.0 ;
# === END ===
END CUT12

LAYER MET2
  TYPE ROUTING ;
  PITCH 0.200 ;
  OFFSET 0.200 ;
  WIDTH 0.100 ;
  MAXWIDTH 3.000 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_MINSTEP "MINSTEP 0.045 MAXEDGES 1 ;" ;
# === END ===
  AREA 0.038 ;
  PROPERTY LEF58_VOLTAGESPACING "VOLTAGESPACING 0.9 0.1 5.0 0.3 ; VOLTAGESPACING TOCUT BELOW 0.9 0.1 5.0 0.5 ; VOLTAGESPACING TOCUT ABOVE 0.9 0.1 5.0 0.5 ;" ;
  MINENCLOSEDAREA 0.110 ;
  MINENCLOSEDAREA 0.800 WIDTH 0.210 ;
  MINENCLOSEDAREA 3.200 WIDTH 1.500 ;
  MINIMUMCUT 2 WIDTH 0.299 ;
  MINIMUMCUT 3 WIDTH 0.699 ;
  MINIMUMCUT 2 WIDTH 0.299 LENGTH 0.774 WITHIN 20000 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.000  0.180  0.380
    WIDTH 0.000        0.100  0.100  0.100
    WIDTH 0.150        0.100  0.120  0.120
    WIDTH 0.180        0.120  0.120  0.120
    WIDTH 0.210        0.120  0.120  0.150
    WIDTH 0.320        0.140  0.140  0.150
    WIDTH 1.500        0.140  0.140  0.500 ;
  MINIMUMDENSITY 20.000 ;
  MAXIMUMDENSITY 80.000 ;
  DENSITYCHECKWINDOW 40.000 40.000 ;
  DENSITYCHECKSTEP 10.000 ;
  DIRECTION VERTICAL ;
# === LEF v5.5 SPEC ===
#  ANTENNACUMAREARATIO 400.0 ;
#  ANTENNACUMDIFFAREARATIO PWL
#   ( ( 0.00000  400.0 ) ( 0.01919 400.0 ) ( 0.01920 100000.000 )
#     ( 1000.00000 100000.000 ) ) ;
#  ANTENNAAREAFACTOR 1.1 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_ANTENNACUMROUTINGPLUSCUT "ANTENNACUMROUTINGPLUSCUT ;" ;
  PROPERTY LEF57_ANTENNAAREAMINUSDIFF "ANTENNAAREAMINUSDIFF 118750 ;" ;
  ANTENNACUMDIFFAREARATIO 2000.0 ;
  ANTENNAAREAFACTOR 1.0 ;
# === END ===
END MET2

LAYER CUT23
  TYPE CUT ;
  SPACING 0.100 ;
# === LEF v5.6 SPEC ===
  ENCLOSURE 0.000 0.040 ;
  ENCLOSURE 0.015 0.040 WIDTH 0.801 ;
  ENCLOSURE 0.035 0.040 WIDTH 1.201 ;
# === END ===
# === LEF v5.5 SPEC ===
#  ANTENNACUMAREARATIO 1600.0 ;
#  ANTENNACUMDIFFAREARATIO PWL
#   ( ( 0.00000  1600.0 ) ( 0.01919 1600.0 ) ( 0.01920 100000.000 )
#     ( 1000.00000 100000.000 ) ) ;
#  ANTENNAAREAFACTOR 100.0 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_ANTENNACUMROUTINGPLUSCUT "ANTENNACUMROUTINGPLUSCUT ;" ;
  PROPERTY LEF57_ANTENNAAREAMINUSDIFF "ANTENNAAREAMINUSDIFF 118750 ;" ;
  ANTENNACUMDIFFAREARATIO 2000.0 ;
  ANTENNAAREAFACTOR 100.0 ;
# === END ===
END CUT23

LAYER MET3
  TYPE ROUTING ;
  PITCH 0.200 ;
  OFFSET 0.200 ;
  WIDTH 0.100 ;
  MAXWIDTH 3.000 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_MINSTEP "MINSTEP 0.045 MAXEDGES 1 ;" ;
# === END ===
  AREA 0.038 ;
  MINENCLOSEDAREA 0.110 ;
  MINENCLOSEDAREA 0.800 WIDTH 0.210 ;
  MINENCLOSEDAREA 3.200 WIDTH 1.500 ;
  MINIMUMCUT 2 WIDTH 0.299 ;
  MINIMUMCUT 3 WIDTH 0.699 ;
  MINIMUMCUT 2 WIDTH 0.299 LENGTH 0.774 WITHIN 20000 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.000  0.180  0.380
    WIDTH 0.000        0.100  0.100  0.100
    WIDTH 0.150        0.100  0.120  0.120
    WIDTH 0.180        0.120  0.120  0.120
    WIDTH 0.210        0.120  0.120  0.150
    WIDTH 0.320        0.140  0.140  0.150
    WIDTH 1.500        0.140  0.140  0.500 ;
  MINIMUMDENSITY 20.000 ;
  MAXIMUMDENSITY 80.000 ;
  DENSITYCHECKWINDOW 40.000 40.000 ;
  DENSITYCHECKSTEP 10.000 ;
  DIRECTION HORIZONTAL ;
# === LEF v5.5 SPEC ===
#  ANTENNACUMAREARATIO 400.0 ;
#  ANTENNACUMDIFFAREARATIO PWL
#   ( ( 0.00000  400.0 ) ( 0.01919 400.0 ) ( 0.01920 100000.000 )
#     ( 1000.00000 100000.000 ) ) ;
#  ANTENNAAREAFACTOR 1.1 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_ANTENNACUMROUTINGPLUSCUT "ANTENNACUMROUTINGPLUSCUT ;" ;
  PROPERTY LEF57_ANTENNAAREAMINUSDIFF "ANTENNAAREAMINUSDIFF 118750 ;" ;
  ANTENNACUMDIFFAREARATIO 2000.0 ;
  ANTENNAAREAFACTOR 1.0 ;
# === END ===
END MET3

LAYER CUT34
  TYPE CUT ;
  SPACING 0.100 ;
# === LEF v5.6 SPEC ===
  ENCLOSURE 0.000 0.040 ;
  ENCLOSURE 0.015 0.040 WIDTH 0.801 ;
  ENCLOSURE 0.035 0.040 WIDTH 1.201 ;
# === END ===
# === LEF v5.5 SPEC ===
#  ANTENNACUMAREARATIO 1600.0 ;
#  ANTENNACUMDIFFAREARATIO PWL
#   ( ( 0.00000  1600.0 ) ( 0.01919 1600.0 ) ( 0.01920 100000.000 )
#     ( 1000.00000 100000.000 ) ) ;
#  ANTENNAAREAFACTOR 100.0 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_ANTENNACUMROUTINGPLUSCUT "ANTENNACUMROUTINGPLUSCUT ;" ;
  PROPERTY LEF57_ANTENNAAREAMINUSDIFF "ANTENNAAREAMINUSDIFF 118750 ;" ;
  ANTENNACUMDIFFAREARATIO 2000.0 ;
  ANTENNAAREAFACTOR 100.0 ;
# === END ===
END CUT34

LAYER MET4
  TYPE ROUTING ;
  PITCH 0.200 ;
  OFFSET 0.200 ;
  WIDTH 0.100 ;
  MAXWIDTH 3.000 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_MINSTEP "MINSTEP 0.045 MAXEDGES 1 ;" ;
# === END ===
  AREA 0.038 ;
  MINENCLOSEDAREA 0.110 ;
  MINENCLOSEDAREA 0.800 WIDTH 0.210 ;
  MINENCLOSEDAREA 3.200 WIDTH 1.500 ;
  MINIMUMCUT 2 WIDTH 0.299 ;
  MINIMUMCUT 3 WIDTH 0.699 ;
  MINIMUMCUT 2 WIDTH 0.299 LENGTH 0.774 WITHIN 20000 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.000  0.180  0.380
    WIDTH 0.000        0.100  0.100  0.100
    WIDTH 0.150        0.100  0.120  0.120
    WIDTH 0.180        0.120  0.120  0.120
    WIDTH 0.210        0.120  0.120  0.150
    WIDTH 0.320        0.140  0.140  0.150
    WIDTH 1.500        0.140  0.140  0.500 ;
  MINIMUMDENSITY 20.000 ;
  MAXIMUMDENSITY 80.000 ;
  DENSITYCHECKWINDOW 40.000 40.000 ;
  DENSITYCHECKSTEP 10.000 ;
  DIRECTION VERTICAL ;
# === LEF v5.5 SPEC ===
#  ANTENNACUMAREARATIO 400.0 ;
#  ANTENNACUMDIFFAREARATIO PWL
#   ( ( 0.00000  400.0 ) ( 0.01919 400.0 ) ( 0.01920 100000.000 )
#     ( 1000.00000 100000.000 ) ) ;
#  ANTENNAAREAFACTOR 1.1 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_ANTENNACUMROUTINGPLUSCUT "ANTENNACUMROUTINGPLUSCUT ;" ;
  PROPERTY LEF57_ANTENNAAREAMINUSDIFF "ANTENNAAREAMINUSDIFF 118750 ;" ;
  ANTENNACUMDIFFAREARATIO 2000.0 ;
  ANTENNAAREAFACTOR 1.0 ;
# === END ===
END MET4

LAYER CUT45
  TYPE CUT ;
  SPACING 0.100 ;
# === LEF v5.6 SPEC ===
  ENCLOSURE 0.000 0.040 ;
  ENCLOSURE 0.015 0.040 WIDTH 0.801 ;
  ENCLOSURE 0.035 0.040 WIDTH 1.201 ;
# === END ===
# === LEF v5.5 SPEC ===
#  ANTENNACUMAREARATIO 1600.0 ;
#  ANTENNACUMDIFFAREARATIO PWL
#   ( ( 0.00000  1600.0 ) ( 0.01919 1600.0 ) ( 0.01920 100000.000 )
#     ( 1000.00000 100000.000 ) ) ;
#  ANTENNAAREAFACTOR 100.0 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_ANTENNACUMROUTINGPLUSCUT "ANTENNACUMROUTINGPLUSCUT ;" ;
  PROPERTY LEF57_ANTENNAAREAMINUSDIFF "ANTENNAAREAMINUSDIFF 118750 ;" ;
  ANTENNACUMDIFFAREARATIO 2000.0 ;
  ANTENNAAREAFACTOR 100.0 ;
# === END ===
END CUT45

LAYER MET5
  TYPE ROUTING ;
  PITCH 0.200 ;
  OFFSET 0.200 ;
  WIDTH 0.100 ;
  MAXWIDTH 3.000 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_MINSTEP "MINSTEP 0.045 MAXEDGES 1 ;" ;
# === END ===
  AREA 0.038 ;
  MINENCLOSEDAREA 0.110 ;
  MINENCLOSEDAREA 0.800 WIDTH 0.210 ;
  MINENCLOSEDAREA 3.200 WIDTH 1.500 ;
  MINIMUMCUT 2 WIDTH 0.299 FROMBELOW ;
  MINIMUMCUT 3 WIDTH 0.699 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 0.299 FROMBELOW LENGTH 0.774 WITHIN 20000 ;
  MINIMUMCUT 2 WIDTH 1.199 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 1.199 FROMABOVE LENGTH 1.199 WITHIN 5.001 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.000  0.180  0.380
    WIDTH 0.000        0.100  0.100  0.100
    WIDTH 0.150        0.100  0.120  0.120
    WIDTH 0.180        0.120  0.120  0.120
    WIDTH 0.210        0.120  0.120  0.150
    WIDTH 0.320        0.140  0.140  0.150
    WIDTH 1.500        0.140  0.140  0.500 ;
  MINIMUMDENSITY 20.000 ;
  MAXIMUMDENSITY 80.000 ;
  DENSITYCHECKWINDOW 40.000 40.000 ;
  DENSITYCHECKSTEP 10.000 ;
  DIRECTION HORIZONTAL ;
# === LEF v5.5 SPEC ===
#  ANTENNACUMAREARATIO 400.0 ;
#  ANTENNACUMDIFFAREARATIO PWL
#   ( ( 0.00000  400.0 ) ( 0.01919 400.0 ) ( 0.01920 100000.000 )
#     ( 1000.00000 100000.000 ) ) ;
#  ANTENNAAREAFACTOR 1.1 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_ANTENNACUMROUTINGPLUSCUT "ANTENNACUMROUTINGPLUSCUT ;" ;
  PROPERTY LEF57_ANTENNAAREAMINUSDIFF "ANTENNAAREAMINUSDIFF 118750 ;" ;
  ANTENNACUMDIFFAREARATIO 2000.0 ;
  ANTENNAAREAFACTOR 1.0 ;
# === END ===
END MET5

LAYER CUTG1
  TYPE CUT ;
  SPACING 0.400 ;
# === LEF v5.6 SPEC ===
  ENCLOSURE BELOW 0.060 0.060 ;
  ENCLOSURE BELOW 0.100 0.100 WIDTH 1.261 ;
  ENCLOSURE ABOVE 0.000 0.000 ;
  ENCLOSURE ABOVE 0.100 0.100 WIDTH 1.401 ;
# === END ===
# === LEF v5.5 SPEC ===
#  ANTENNACUMAREARATIO 1600.0 ;
#  ANTENNACUMDIFFAREARATIO PWL
#   ( ( 0.00000  1600.0 ) ( 0.01919 1600.0 ) ( 0.01920 100000.000 )
#     ( 1000.00000 100000.000 ) ) ;
#  ANTENNAAREAFACTOR 7.5 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_ANTENNACUMROUTINGPLUSCUT "ANTENNACUMROUTINGPLUSCUT ;" ;
  PROPERTY LEF57_ANTENNAAREAMINUSDIFF "ANTENNAAREAMINUSDIFF 118750 ;" ;
  ANTENNACUMDIFFAREARATIO 2000.0 ;
  ANTENNAAREAFACTOR 7.5 ;
# === END ===
END CUTG1

LAYER METG1
  TYPE ROUTING ;
  PITCH 0.800 ;
  OFFSET 0.200 ;
  WIDTH 0.400 ;
  MAXWIDTH 12.000 ;
  AREA 0.480 ;
  MINENCLOSEDAREA 2.800 ;
  MINENCLOSEDAREA 16.000 WIDTH 1.600 ;
  MINENCLOSEDAREA 36.000 WIDTH 4.600 ;
  MINENCLOSEDAREA 100.000 WIDTH 6.000 ;
  MINENCLOSEDAREA 225.000 WIDTH 10.000 ;
  MINIMUMCUT 2 WIDTH 1.199 FROMBELOW ;
  MINIMUMCUT 2 WIDTH 1.199 FROMBELOW LENGTH 1.199 WITHIN 5.001 ;
  MINIMUMCUT 2 WIDTH 2.399 FROMABOVE ;
  MINIMUMCUT 2 WIDTH 2.399 FROMABOVE LENGTH 2.399 WITHIN 5.001 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.000  100.0
    WIDTH 0.000        0.400  0.400
    WIDTH 1.600        0.500  0.500
    WIDTH 4.600        0.900  0.900
    WIDTH 6.000        2.500  2.500
    WIDTH 10.00        3.750  3.750 ;
  MINIMUMDENSITY 20.000 ;
  MAXIMUMDENSITY 80.000 ;
  DENSITYCHECKWINDOW 40.000 40.000 ;
  DENSITYCHECKSTEP 10.000 ;
  DIRECTION VERTICAL ;
# === LEF v5.5 SPEC ===
#  ANTENNACUMAREARATIO 400.0 ;
#  ANTENNACUMDIFFAREARATIO PWL
#   ( ( 0.00000  400.0 ) ( 0.01919 400.0 ) ( 0.01920 100000.000 )
#     ( 1000.00000 100000.000 ) ) ;
#  ANTENNAAREAFACTOR 1.1 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_ANTENNACUMROUTINGPLUSCUT "ANTENNACUMROUTINGPLUSCUT ;" ;
  PROPERTY LEF57_ANTENNAAREAMINUSDIFF "ANTENNAAREAMINUSDIFF 118750 ;" ;
  ANTENNACUMDIFFAREARATIO 2000.0 ;
  ANTENNAAREAFACTOR 1.0 ;
# === END ===
END METG1

LAYER CUTTOP
  TYPE CUT ;
  SPACING 1.100 ;
# === LEF v5.6 SPEC === 
  ENCLOSURE BELOW 0.100 0.100 ;
  ENCLOSURE ABOVE 0.250 0.250 ;
# === END ===
# === LEF v5.5 SPEC ===
#  ANTENNACUMAREARATIO 1600.0 ;
#  ANTENNACUMDIFFAREARATIO PWL
#   ( ( 0.00000  1600.0 ) ( 0.01919 1600.0 ) ( 0.01920 100000.000 )
#     ( 1000.00000 100000.000 ) ) ;
#  ANTENNAAREAFACTOR 12.0 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_ANTENNACUMROUTINGPLUSCUT "ANTENNACUMROUTINGPLUSCUT ;" ;
  PROPERTY LEF57_ANTENNAAREAMINUSDIFF "ANTENNAAREAMINUSDIFF 118750 ;" ;
  ANTENNACUMDIFFAREARATIO 2000.0 ;
  ANTENNAAREAFACTOR 12.0 ;
# === END ===
END CUTTOP

LAYER METTOP
  TYPE ROUTING ;
  PITCH 1.600 ;
  OFFSET 0.200 ;
  WIDTH 0.800 ;
  MAXWIDTH 30.000 ;
  AREA 1.890 ;
  MINENCLOSEDAREA 4.000 ;
#  MINIMUMCUT 2 WIDTH 2.399 ;
#  MINIMUMCUT 2 WIDTH 2.399 LENGTH 2.399 WITHIN 5.001 ;
  SPACINGTABLE
    PARALLELRUNLENGTH  0.000  100.0
    WIDTH  0.000       0.800  0.800
    WIDTH 99.999       1.120  1.120 ;
  MINIMUMDENSITY 30.000 ;
  MAXIMUMDENSITY 85.000 ;
  DIRECTION HORIZONTAL ;
# === LEF v5.5 SPEC ===
#  ANTENNACUMAREARATIO 400.0 ;
#  ANTENNACUMDIFFAREARATIO PWL
#   ( ( 0.00000  400.0 ) ( 0.01919 400.0 ) ( 0.01920 100000.000 )
#     ( 1000.00000 100000.000 ) ) ;
#  ANTENNAAREAFACTOR 1.1 ;
# === LEF v5.6 SPEC ===
  PROPERTY LEF57_ANTENNACUMROUTINGPLUSCUT "ANTENNACUMROUTINGPLUSCUT ;" ;
  PROPERTY LEF57_ANTENNAAREAMINUSDIFF "ANTENNAAREAMINUSDIFF 118750 ;" ;
  ANTENNACUMDIFFAREARATIO 2000.0 ;
  ANTENNAAREAFACTOR 1.0 ;
# === END ===
END METTOP

LAYER OVLAP
  TYPE OVERLAP ;
END OVLAP

# POWER-RAIL VIA
VIA VIA34P
  LAYER MET3 ;
    RECT -0.725 -0.150  0.725  0.150 ;
  LAYER CUT34 ;
    RECT -0.650 -0.150 -0.550 -0.050 ;
    RECT -0.450 -0.150 -0.350 -0.050 ;
    RECT -0.250 -0.150 -0.150 -0.050 ;
    RECT -0.050 -0.150  0.050 -0.050 ;
    RECT  0.150 -0.150  0.250 -0.050 ;
    RECT  0.350 -0.150  0.450 -0.050 ;
    RECT  0.550 -0.150  0.650 -0.050 ;
    RECT -0.650  0.050 -0.550  0.150 ;
    RECT -0.450  0.050 -0.350  0.150 ;
    RECT -0.250  0.050 -0.150  0.150 ;
    RECT -0.050  0.050  0.050  0.150 ;
    RECT  0.150  0.050  0.250  0.150 ;
    RECT  0.350  0.050  0.450  0.150 ;
    RECT  0.550  0.050  0.650  0.150 ;
  LAYER MET4 ;
    RECT -0.725 -0.185  0.725  0.185 ;
END VIA34P

VIA VIA34P2
  LAYER MET3 ;
    RECT -0.725 -0.160  0.725  0.160 ;
  LAYER CUT34 ;
    RECT -0.650 -0.150 -0.550 -0.050 ;
    RECT -0.450 -0.150 -0.350 -0.050 ;
    RECT -0.250 -0.150 -0.150 -0.050 ;
    RECT -0.050 -0.150  0.050 -0.050 ;
    RECT  0.150 -0.150  0.250 -0.050 ;
    RECT  0.350 -0.150  0.450 -0.050 ;
    RECT  0.550 -0.150  0.650 -0.050 ;
    RECT -0.650  0.050 -0.550  0.150 ;
    RECT -0.450  0.050 -0.350  0.150 ;
    RECT -0.250  0.050 -0.150  0.150 ;
    RECT -0.050  0.050  0.050  0.150 ;
    RECT  0.150  0.050  0.250  0.150 ;
    RECT  0.350  0.050  0.450  0.150 ;
    RECT  0.550  0.050  0.650  0.150 ;
  LAYER MET4 ;
    RECT -0.725 -0.185  0.725  0.185 ;
END VIA34P2

# SINGLE-VIA
VIA VIA1_HV DEFAULT
  LAYER MET1 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA1_HV

VIA VIA1_HH DEFAULT
  LAYER MET1 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA1_HH

VIA VIA1_VH DEFAULT
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA1_VH

VIA VIA1_VV DEFAULT
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA1_VV

# MULTI-VIA
VIA VIA1_2N DEFAULT
  LAYER MET1 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA1_2N

VIA VIA1_2NV DEFAULT
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA1_2NV

VIA VIA1_2NR DEFAULT
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA1_2NR

VIA VIA1_2S DEFAULT
  LAYER MET1 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA1_2S

VIA VIA1_2SV DEFAULT
  LAYER MET1 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA1_2SV

VIA VIA1_2SR DEFAULT
  LAYER MET1 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA1_2SR

VIA VIA1_2V DEFAULT
  LAYER MET1 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA1_2V

VIA VIA1_2CV DEFAULT
  LAYER MET1 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA1_2CV

VIA VIA1_2VR DEFAULT
  LAYER MET1 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA1_2VR

VIA VIA1_2E DEFAULT
  LAYER MET1 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA1_2E

VIA VIA1_2EH DEFAULT
  LAYER MET1 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA1_2EH

VIA VIA1_2ER DEFAULT
  LAYER MET1 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA1_2ER

VIA VIA1_2W DEFAULT
  LAYER MET1 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA1_2W

VIA VIA1_2WH DEFAULT
  LAYER MET1 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA1_2WH

VIA VIA1_2WR DEFAULT
  LAYER MET1 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA1_2WR

VIA VIA1_2H DEFAULT
  LAYER MET1 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA1_2H

VIA VIA1_2CH DEFAULT
  LAYER MET1 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA1_2CH

VIA VIA1_2HR DEFAULT
  LAYER MET1 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA1_2HR

VIA VIA1_3H DEFAULT
  LAYER MET1 ;
    RECT -0.290 -0.050  0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.250 -0.090  0.250 0.090 ;
END VIA1_3H

VIA VIA1_3V DEFAULT
  LAYER MET1 ;
    RECT -0.090 -0.250 0.090  0.250 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.290 ;
END VIA1_3V

VIA VIA1_4H DEFAULT
  LAYER MET1 ;
    RECT -0.390 -0.050  0.390 0.050 ;
  LAYER CUT12 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET2 ;
    RECT -0.350 -0.090  0.350 0.090 ;
END VIA1_4H

VIA VIA1_4V DEFAULT
  LAYER MET1 ;
    RECT -0.090 -0.350 0.090  0.350 ;
  LAYER CUT12 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET2 ;
    RECT -0.050 -0.390 0.050  0.390 ;
END VIA1_4V

# SINGLE-VIA
VIA VIA2_VH DEFAULT
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA2_VH

VIA VIA2_VV DEFAULT
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA2_VV

VIA VIA2_HV DEFAULT
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA2_HV

VIA VIA2_HH DEFAULT
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA2_HH

# STACK-VIA
VIA VIA2_NS DEFAULT
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA2_NS

VIA VIA2_SS DEFAULT
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050 0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA2_SS

VIA VIA2_VS DEFAULT
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050 0.190 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA2_VS

# MULTI-VIA
VIA VIA2_2N DEFAULT
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA2_2N

VIA VIA2_2S DEFAULT
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA2_2S

VIA VIA2_2V DEFAULT
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA2_2V

VIA VIA2_2E DEFAULT
  LAYER MET2 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA2_2E

VIA VIA2_2W DEFAULT
  LAYER MET2 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA2_2W

VIA VIA2_2H DEFAULT
  LAYER MET2 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA2_2H

VIA VIA2_2NR DEFAULT
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA2_2NR

VIA VIA2_2SR DEFAULT
  LAYER MET2 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA2_2SR

VIA VIA2_2VR DEFAULT
  LAYER MET2 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA2_2VR

VIA VIA2_2ER DEFAULT
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA2_2ER

VIA VIA2_2WR DEFAULT
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA2_2WR

VIA VIA2_2HR DEFAULT
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA2_2HR

VIA VIA2_2NV DEFAULT
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA2_2NV

VIA VIA2_2SV DEFAULT
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA2_2SV

VIA VIA2_2CV DEFAULT
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA2_2CV

VIA VIA2_2EH DEFAULT
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA2_2EH

VIA VIA2_2WH DEFAULT
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA2_2WH

VIA VIA2_2CH DEFAULT
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA2_2CH

VIA VIA2_3H DEFAULT
  LAYER MET2 ;
    RECT -0.250 -0.090  0.250 0.090 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.290 0.050 ;
END VIA2_3H

VIA VIA2_3V DEFAULT
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.250 ;
END VIA2_3V

VIA VIA2_4H DEFAULT
  LAYER MET2 ;
    RECT -0.350 -0.090  0.350 0.090 ;
  LAYER CUT23 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET3 ;
    RECT -0.390 -0.050  0.390 0.050 ;
END VIA2_4H

VIA VIA2_4V DEFAULT
  LAYER MET2 ;
    RECT -0.050 -0.390 0.050  0.390 ;
  LAYER CUT23 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET3 ;
    RECT -0.090 -0.350 0.090  0.350 ;
END VIA2_4V

# SINGLE-VIA
VIA VIA3_HV DEFAULT
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA3_HV

VIA VIA3_HH DEFAULT
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA3_HH

VIA VIA3_VH DEFAULT
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA3_VH

VIA VIA3_VV DEFAULT
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA3_VV

# STACK-VIA
VIA VIA3_ES DEFAULT
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA3_ES

VIA VIA3_WS DEFAULT
  LAYER MET3 ;
    RECT -0.290 -0.050 0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA3_WS

VIA VIA3_HS DEFAULT
  LAYER MET3 ;
    RECT -0.190 -0.050 0.190 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA3_HS

# MULTI-VIA
VIA VIA3_2N DEFAULT
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA3_2N

VIA VIA3_2S DEFAULT
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA3_2S

VIA VIA3_2V DEFAULT
  LAYER MET3 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT34 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA3_2V

VIA VIA3_2E DEFAULT
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA3_2E

VIA VIA3_2W DEFAULT
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA3_2W

VIA VIA3_2H DEFAULT
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT34 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET4 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA3_2H

VIA VIA3_2NR DEFAULT
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA3_2NR

VIA VIA3_2SR DEFAULT
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA3_2SR

VIA VIA3_2VR DEFAULT
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT34 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET4 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA3_2VR

VIA VIA3_2ER DEFAULT
  LAYER MET3 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA3_2ER

VIA VIA3_2WR DEFAULT
  LAYER MET3 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA3_2WR

VIA VIA3_2HR DEFAULT
  LAYER MET3 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT34 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET4 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA3_2HR

VIA VIA3_2NV DEFAULT
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA3_2NV

VIA VIA3_2SV DEFAULT
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA3_2SV

VIA VIA3_2CV DEFAULT
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT34 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA3_2CV

VIA VIA3_2EH DEFAULT
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA3_2EH

VIA VIA3_2WH DEFAULT
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA3_2WH

VIA VIA3_2CH DEFAULT
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT34 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET4 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA3_2CH

VIA VIA3_3H DEFAULT
  LAYER MET3 ;
    RECT -0.290 -0.050  0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.250 -0.090  0.250 0.090 ;
END VIA3_3H

VIA VIA3_3V DEFAULT
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.250 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.290 ;
END VIA3_3V

VIA VIA3_4H DEFAULT
  LAYER MET3 ;
    RECT -0.390 -0.050  0.390 0.050 ;
  LAYER CUT34 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET4 ;
    RECT -0.350 -0.090  0.350 0.090 ;
END VIA3_4H

VIA VIA3_4V DEFAULT
  LAYER MET3 ;
    RECT -0.090 -0.350 0.090  0.350 ;
  LAYER CUT34 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET4 ;
    RECT -0.050 -0.390 0.050  0.390 ;
END VIA3_4V

# SINGLE-VIA
VIA VIA4_VH DEFAULT
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA4_VH

VIA VIA4_VV DEFAULT
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA4_VV

VIA VIA4_HV DEFAULT
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA4_HV

VIA VIA4_HH DEFAULT
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA4_HH

# STACK-VIA
VIA VIA4_NS DEFAULT
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA4_NS

VIA VIA4_SS DEFAULT
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050 0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA4_SS

VIA VIA4_VS DEFAULT
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050 0.190 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA4_VS

# MULTI-VIA
VIA VIA4_2N DEFAULT
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA4_2N

VIA VIA4_2S DEFAULT
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA4_2S

VIA VIA4_2V DEFAULT
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT45 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET5 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA4_2V

VIA VIA4_2E DEFAULT
  LAYER MET4 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA4_2E

VIA VIA4_2W DEFAULT
  LAYER MET4 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA4_2W

VIA VIA4_2H DEFAULT
  LAYER MET4 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT45 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET5 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA4_2H

VIA VIA4_2NR DEFAULT
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA4_2NR

VIA VIA4_2SR DEFAULT
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA4_2SR

VIA VIA4_2VR DEFAULT
  LAYER MET4 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT45 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET5 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA4_2VR

VIA VIA4_2ER DEFAULT
  LAYER MET4 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA4_2ER

VIA VIA4_2WR DEFAULT
  LAYER MET4 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA4_2WR

VIA VIA4_2HR DEFAULT
  LAYER MET4 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT45 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET5 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA4_2HR

VIA VIA4_2NV DEFAULT
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA4_2NV

VIA VIA4_2SV DEFAULT
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA4_2SV

VIA VIA4_2CV DEFAULT
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT45 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET5 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA4_2CV

VIA VIA4_2EH DEFAULT
  LAYER MET4 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA4_2EH

VIA VIA4_2WH DEFAULT
  LAYER MET4 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA4_2WH

VIA VIA4_2CH DEFAULT
  LAYER MET4 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT45 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET5 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA4_2CH

VIA VIA4_3H DEFAULT
  LAYER MET4 ;
    RECT -0.250 -0.090  0.250 0.090 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.290 -0.050  0.290 0.050 ;
END VIA4_3H

VIA VIA4_3V DEFAULT
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.290 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET5 ;
    RECT -0.090 -0.250 0.090  0.250 ;
END VIA4_3V

VIA VIA4_4H DEFAULT
  LAYER MET4 ;
    RECT -0.350 -0.090  0.350 0.090 ;
  LAYER CUT45 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET5 ;
    RECT -0.390 -0.050  0.390 0.050 ;
END VIA4_4H

VIA VIA4_4V DEFAULT
  LAYER MET4 ;
    RECT -0.050 -0.390 0.050  0.390 ;
  LAYER CUT45 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET5 ;
    RECT -0.090 -0.350 0.090  0.350 ;
END VIA4_4V

# SINGLE/STACK-VIA
VIA VIAG1 DEFAULT
  LAYER MET5 ;
    RECT -0.260 -0.260 0.260 0.260 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER METG1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
END VIAG1

VIA VIAG1_N DEFAULT
  LAYER MET5 ;
    RECT -0.260 -0.200 0.260 0.320 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.140 0.200 0.260 ;
  LAYER METG1 ;
    RECT -0.200 -0.140 0.200 0.260 ;
END VIAG1_N

VIA VIAG1_S DEFAULT
  LAYER MET5 ;
    RECT -0.260 -0.320 0.260 0.200 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.260 0.200 0.140 ;
  LAYER METG1 ;
    RECT -0.200 -0.260 0.200 0.140 ;
END VIAG1_S

VIA VIAG1_E DEFAULT
  LAYER MET5 ;
    RECT -0.200 -0.260 0.320 0.260 ;
  LAYER CUTG1 ;
    RECT -0.140 -0.200 0.260 0.200 ;
  LAYER METG1 ;
    RECT -0.140 -0.200 0.260 0.200 ;
END VIAG1_E

VIA VIAG1_W DEFAULT
  LAYER MET5 ;
    RECT -0.320 -0.260 0.200 0.260 ;
  LAYER CUTG1 ;
    RECT -0.260 -0.200 0.140 0.200 ;
  LAYER METG1 ;
    RECT -0.260 -0.200 0.140 0.200 ;
END VIAG1_W

# MULTI-VIA
VIA VIAG1_2N DEFAULT
  LAYER MET5 ;
    RECT -0.260 -0.260 0.260 1.060 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
    RECT -0.200  0.600 0.200 1.000 ;
  LAYER METG1 ;
    RECT -0.200 -0.200 0.200 1.000 ;
END VIAG1_2N

VIA VIAG1_2S DEFAULT
  LAYER MET5 ;
    RECT -0.260 -1.060 0.260  0.260 ;
  LAYER CUTG1 ;
    RECT -0.200 -1.000 0.200 -0.600 ;
    RECT -0.200 -0.200 0.200  0.200 ;
  LAYER METG1 ;
    RECT -0.200 -1.000 0.200  0.200 ;
END VIAG1_2S

VIA VIAG1_2V DEFAULT
  LAYER MET5 ;
    RECT -0.260 -0.660 0.260  0.660 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.600 0.200 -0.200 ;
    RECT -0.200  0.200 0.200  0.600 ;
  LAYER METG1 ;
    RECT -0.200 -0.600 0.200  0.600 ;
END VIAG1_2V

VIA VIAG1_2E DEFAULT
  LAYER MET5 ;
    RECT -0.260 -0.260 1.060  0.260 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200  0.200 ;
    RECT  0.600 -0.200 1.000  0.200 ;
  LAYER METG1 ;
    RECT -0.200 -0.200 1.000  0.200 ;
END VIAG1_2E

VIA VIAG1_2W DEFAULT
  LAYER MET5 ;
    RECT -1.060 -0.260  0.260 0.260 ;
  LAYER CUTG1 ;
    RECT -1.000 -0.200 -0.600 0.200 ;
    RECT -0.200 -0.200  0.200 0.200 ;
  LAYER METG1 ;
    RECT -1.000 -0.200  0.200 0.200 ;
END VIAG1_2W

VIA VIAG1_2H DEFAULT
  LAYER MET5 ;
    RECT -0.660 -0.260  0.660 0.260 ;
  LAYER CUTG1 ;
    RECT -0.600 -0.200 -0.200 0.200 ;
    RECT  0.200 -0.200  0.600 0.200 ;
  LAYER METG1 ;
    RECT -0.600 -0.200  0.600 0.200 ;
END VIAG1_2H

# SINGLE/STACK-VIA
VIA VIATOP DEFAULT
  LAYER METG1 ;
    RECT -0.350 -0.350 0.350 0.350 ;
  LAYER CUTTOP ;
    RECT -0.250 -0.250 0.250 0.250 ;
  LAYER METTOP ;
    RECT -0.500 -0.500 0.500 0.500 ;
END VIATOP

# MULTI-VIA
VIA VIATOP_2N DEFAULT
  LAYER METG1 ;
    RECT -0.350 -0.350 0.350 1.950 ;
  LAYER CUTTOP ;
    RECT -0.250 -0.250 0.250 0.250 ;
    RECT -0.250  1.350 0.250 1.850 ;
  LAYER METTOP ;
    RECT -0.500 -0.500 0.500 2.100 ;
END VIATOP_2N

VIA VIATOP_2S DEFAULT
  LAYER METG1 ;
    RECT -0.350 -1.950 0.350  0.350 ;
  LAYER CUTTOP ;
    RECT -0.250 -1.850 0.250 -1.350 ;
    RECT -0.250 -0.250 0.250  0.250 ;
  LAYER METTOP ;
    RECT -0.500 -2.100 0.500  0.500 ;
END VIATOP_2S

VIA VIATOP_2V DEFAULT
  LAYER METG1 ;
    RECT -0.350 -1.150 0.350  1.150 ;
  LAYER CUTTOP ;
    RECT -0.250 -1.050 0.250 -0.550 ;
    RECT -0.250  0.550 0.250  1.050 ;
  LAYER METTOP ;
    RECT -0.500 -1.300 0.500  1.300 ;
END VIATOP_2V

VIA VIATOP_2E DEFAULT
  LAYER METG1 ;
    RECT -0.350 -0.350 1.950 0.350 ;
  LAYER CUTTOP ;
    RECT -0.250 -0.250 0.250 0.250 ;
    RECT  1.350 -0.250 1.850 0.250 ;
  LAYER METTOP ;
    RECT -0.500 -0.500 2.100 0.500 ;
END VIATOP_2E

VIA VIATOP_2W DEFAULT
  LAYER METG1 ;
    RECT -1.950 -0.350  0.350 0.350 ;
  LAYER CUTTOP ;
    RECT -1.850 -0.250 -1.350 0.250 ;
    RECT -0.250 -0.250  0.250 0.250 ;
  LAYER METTOP ;
    RECT -2.100 -0.500  0.500 0.500 ;
END VIATOP_2W

VIA VIATOP_2H DEFAULT
  LAYER METG1 ;
    RECT -1.150 -0.350  1.150 0.350 ;
  LAYER CUTTOP ;
    RECT -1.050 -0.250 -0.550 0.250 ;
    RECT  0.550 -0.250  1.050 0.250 ;
  LAYER METTOP ;
    RECT -1.300 -0.500  1.300 0.500 ;
END VIATOP_2H

SPACING
  SAMENET CUT01 CUT12 0.000 STACK ;
  SAMENET CUT12 CUT23 0.000 STACK ;
  SAMENET CUT23 CUT34 0.000 STACK ;
  SAMENET CUT34 CUT45 0.000 STACK ;
  SAMENET CUT45 CUTG1 0.000 STACK ;
  SAMENET CUTG1 CUTTOP 0.000 STACK ;
END SPACING

NONDEFAULTRULE DOUBLESPACE
LAYER MET1
  WIDTH 0.100 ;
  SPACING 0.200 ;
END MET1

LAYER MET2
  WIDTH 0.100 ;
  SPACING 0.200 ;
END MET2

LAYER MET3
  WIDTH 0.100 ;
  SPACING 0.200 ;
END MET3

LAYER MET4
  WIDTH 0.100 ;
  SPACING 0.200 ;
END MET4

LAYER MET5
  WIDTH 0.100 ;
  SPACING 0.200 ;
END MET5

LAYER METG1
  WIDTH 0.400 ;
  SPACING 0.800 ;
END METG1

LAYER METTOP
  WIDTH 0.800 ;
  SPACING 1.600 ;
END METTOP

# SINGLE-VIA
VIA VIA1_HV_DS
  LAYER MET1 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA1_HV_DS

VIA VIA1_HH_DS
  LAYER MET1 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA1_HH_DS

VIA VIA1_VH_DS
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA1_VH_DS

VIA VIA1_VV_DS
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA1_VV_DS

# MULTI-VIA
VIA VIA1_2N_DS
  LAYER MET1 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA1_2N_DS

VIA VIA1_2NV_DS
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA1_2NV_DS

VIA VIA1_2NR_DS
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA1_2NR_DS

VIA VIA1_2S_DS
  LAYER MET1 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA1_2S_DS

VIA VIA1_2SV_DS
  LAYER MET1 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA1_2SV_DS

VIA VIA1_2SR_DS
  LAYER MET1 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA1_2SR_DS

VIA VIA1_2V_DS
  LAYER MET1 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA1_2V_DS

VIA VIA1_2CV_DS
  LAYER MET1 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA1_2CV_DS

VIA VIA1_2VR_DS
  LAYER MET1 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA1_2VR_DS

VIA VIA1_2E_DS
  LAYER MET1 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA1_2E_DS

VIA VIA1_2EH_DS
  LAYER MET1 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA1_2EH_DS

VIA VIA1_2ER_DS
  LAYER MET1 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA1_2ER_DS

VIA VIA1_2W_DS
  LAYER MET1 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA1_2W_DS

VIA VIA1_2WH_DS
  LAYER MET1 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA1_2WH_DS

VIA VIA1_2WR_DS
  LAYER MET1 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA1_2WR_DS

VIA VIA1_2H_DS
  LAYER MET1 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA1_2H_DS

VIA VIA1_2CH_DS
  LAYER MET1 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA1_2CH_DS

VIA VIA1_2HR_DS
  LAYER MET1 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA1_2HR_DS

VIA VIA1_3H_DS
  LAYER MET1 ;
    RECT -0.290 -0.050  0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.250 -0.090  0.250 0.090 ;
END VIA1_3H_DS

VIA VIA1_3V_DS
  LAYER MET1 ;
    RECT -0.090 -0.250 0.090  0.250 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.290 ;
END VIA1_3V_DS

VIA VIA1_4H_DS
  LAYER MET1 ;
    RECT -0.390 -0.050  0.390 0.050 ;
  LAYER CUT12 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET2 ;
    RECT -0.350 -0.090  0.350 0.090 ;
END VIA1_4H_DS

VIA VIA1_4V_DS
  LAYER MET1 ;
    RECT -0.090 -0.350 0.090  0.350 ;
  LAYER CUT12 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET2 ;
    RECT -0.050 -0.390 0.050  0.390 ;
END VIA1_4V_DS

# SINGLE-VIA
VIA VIA2_VH_DS
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA2_VH_DS

VIA VIA2_VV_DS
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA2_VV_DS

VIA VIA2_HV_DS
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA2_HV_DS

VIA VIA2_HH_DS
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA2_HH_DS

# STACK-VIA
VIA VIA2_NS_DS
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA2_NS_DS

VIA VIA2_SS_DS
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050 0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA2_SS_DS

VIA VIA2_VS_DS
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050 0.190 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA2_VS_DS

# MULTI-VIA
VIA VIA2_2N_DS
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA2_2N_DS

VIA VIA2_2S_DS
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA2_2S_DS

VIA VIA2_2V_DS
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA2_2V_DS

VIA VIA2_2E_DS
  LAYER MET2 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA2_2E_DS

VIA VIA2_2W_DS
  LAYER MET2 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA2_2W_DS

VIA VIA2_2H_DS
  LAYER MET2 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA2_2H_DS

VIA VIA2_2NR_DS
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA2_2NR_DS

VIA VIA2_2SR_DS
  LAYER MET2 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA2_2SR_DS

VIA VIA2_2VR_DS
  LAYER MET2 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA2_2VR_DS

VIA VIA2_2ER_DS
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA2_2ER_DS

VIA VIA2_2WR_DS
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA2_2WR_DS

VIA VIA2_2HR_DS
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA2_2HR_DS

VIA VIA2_2NV_DS
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA2_2NV_DS

VIA VIA2_2SV_DS
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA2_2SV_DS

VIA VIA2_2CV_DS
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA2_2CV_DS

VIA VIA2_2EH_DS
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA2_2EH_DS

VIA VIA2_2WH_DS
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA2_2WH_DS

VIA VIA2_2CH_DS
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA2_2CH_DS

VIA VIA2_3H_DS
  LAYER MET2 ;
    RECT -0.250 -0.090  0.250 0.090 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.290 0.050 ;
END VIA2_3H_DS

VIA VIA2_3V_DS
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.250 ;
END VIA2_3V_DS

VIA VIA2_4H_DS
  LAYER MET2 ;
    RECT -0.350 -0.090  0.350 0.090 ;
  LAYER CUT23 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET3 ;
    RECT -0.390 -0.050  0.390 0.050 ;
END VIA2_4H_DS

VIA VIA2_4V_DS
  LAYER MET2 ;
    RECT -0.050 -0.390 0.050  0.390 ;
  LAYER CUT23 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET3 ;
    RECT -0.090 -0.350 0.090  0.350 ;
END VIA2_4V_DS

# SINGLE-VIA
VIA VIA3_HV_DS
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA3_HV_DS

VIA VIA3_HH_DS
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA3_HH_DS

VIA VIA3_VH_DS
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA3_VH_DS

VIA VIA3_VV_DS
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA3_VV_DS

# STACK-VIA
VIA VIA3_ES_DS
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA3_ES_DS

VIA VIA3_WS_DS
  LAYER MET3 ;
    RECT -0.290 -0.050 0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA3_WS_DS

VIA VIA3_HS_DS
  LAYER MET3 ;
    RECT -0.190 -0.050 0.190 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA3_HS_DS

# MULTI-VIA
VIA VIA3_2N_DS
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA3_2N_DS

VIA VIA3_2S_DS
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA3_2S_DS

VIA VIA3_2V_DS
  LAYER MET3 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT34 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA3_2V_DS

VIA VIA3_2E_DS
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA3_2E_DS

VIA VIA3_2W_DS
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA3_2W_DS

VIA VIA3_2H_DS
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT34 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET4 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA3_2H_DS

VIA VIA3_2NR_DS
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA3_2NR_DS

VIA VIA3_2SR_DS
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA3_2SR_DS

VIA VIA3_2VR_DS
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT34 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET4 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA3_2VR_DS

VIA VIA3_2ER_DS
  LAYER MET3 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA3_2ER_DS

VIA VIA3_2WR_DS
  LAYER MET3 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA3_2WR_DS

VIA VIA3_2HR_DS
  LAYER MET3 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT34 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET4 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA3_2HR_DS

VIA VIA3_2NV_DS
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA3_2NV_DS

VIA VIA3_2SV_DS
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA3_2SV_DS

VIA VIA3_2CV_DS
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT34 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA3_2CV_DS

VIA VIA3_2EH_DS
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA3_2EH_DS

VIA VIA3_2WH_DS
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA3_2WH_DS

VIA VIA3_2CH_DS
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT34 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET4 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA3_2CH_DS

VIA VIA3_3H_DS
  LAYER MET3 ;
    RECT -0.290 -0.050  0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.250 -0.090  0.250 0.090 ;
END VIA3_3H_DS

VIA VIA3_3V_DS
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.250 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.290 ;
END VIA3_3V_DS

VIA VIA3_4H_DS
  LAYER MET3 ;
    RECT -0.390 -0.050  0.390 0.050 ;
  LAYER CUT34 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET4 ;
    RECT -0.350 -0.090  0.350 0.090 ;
END VIA3_4H_DS

VIA VIA3_4V_DS
  LAYER MET3 ;
    RECT -0.090 -0.350 0.090  0.350 ;
  LAYER CUT34 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET4 ;
    RECT -0.050 -0.390 0.050  0.390 ;
END VIA3_4V_DS

# SINGLE-VIA
VIA VIA4_VH_DS
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA4_VH_DS

VIA VIA4_VV_DS
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA4_VV_DS

VIA VIA4_HV_DS
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA4_HV_DS

VIA VIA4_HH_DS
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA4_HH_DS

# STACK-VIA
VIA VIA4_NS_DS
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA4_NS_DS

VIA VIA4_SS_DS
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050 0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA4_SS_DS

VIA VIA4_VS_DS
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050 0.190 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA4_VS_DS

# MULTI-VIA
VIA VIA4_2N_DS
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA4_2N_DS

VIA VIA4_2S_DS
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA4_2S_DS

VIA VIA4_2V_DS
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT45 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET5 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA4_2V_DS

VIA VIA4_2E_DS
  LAYER MET4 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA4_2E_DS

VIA VIA4_2W_DS
  LAYER MET4 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA4_2W_DS

VIA VIA4_2H_DS
  LAYER MET4 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT45 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET5 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA4_2H_DS

VIA VIA4_2NR_DS
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA4_2NR_DS

VIA VIA4_2SR_DS
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA4_2SR_DS

VIA VIA4_2VR_DS
  LAYER MET4 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT45 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET5 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA4_2VR_DS

VIA VIA4_2ER_DS
  LAYER MET4 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA4_2ER_DS

VIA VIA4_2WR_DS
  LAYER MET4 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA4_2WR_DS

VIA VIA4_2HR_DS
  LAYER MET4 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT45 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET5 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA4_2HR_DS

VIA VIA4_2NV_DS
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA4_2NV_DS

VIA VIA4_2SV_DS
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA4_2SV_DS

VIA VIA4_2CV_DS
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT45 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET5 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA4_2CV_DS

VIA VIA4_2EH_DS
  LAYER MET4 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA4_2EH_DS

VIA VIA4_2WH_DS
  LAYER MET4 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA4_2WH_DS

VIA VIA4_2CH_DS
  LAYER MET4 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT45 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET5 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA4_2CH_DS

VIA VIA4_3H_DS
  LAYER MET4 ;
    RECT -0.250 -0.090  0.250 0.090 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.290 -0.050  0.290 0.050 ;
END VIA4_3H_DS

VIA VIA4_3V_DS
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.290 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET5 ;
    RECT -0.090 -0.250 0.090  0.250 ;
END VIA4_3V_DS

VIA VIA4_4H_DS
  LAYER MET4 ;
    RECT -0.350 -0.090  0.350 0.090 ;
  LAYER CUT45 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET5 ;
    RECT -0.390 -0.050  0.390 0.050 ;
END VIA4_4H_DS

VIA VIA4_4V_DS
  LAYER MET4 ;
    RECT -0.050 -0.390 0.050  0.390 ;
  LAYER CUT45 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET5 ;
    RECT -0.090 -0.350 0.090  0.350 ;
END VIA4_4V_DS

# SINGLE/STACK-VIA
VIA VIAG1_DS
  LAYER MET5 ;
    RECT -0.260 -0.260 0.260 0.260 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER METG1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
END VIAG1_DS

VIA VIAG1_N_DS
  LAYER MET5 ;
    RECT -0.260 -0.200 0.260 0.320 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.140 0.200 0.260 ;
  LAYER METG1 ;
    RECT -0.200 -0.140 0.200 0.260 ;
END VIAG1_N_DS

VIA VIAG1_S_DS
  LAYER MET5 ;
    RECT -0.260 -0.320 0.260 0.200 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.260 0.200 0.140 ;
  LAYER METG1 ;
    RECT -0.200 -0.260 0.200 0.140 ;
END VIAG1_S_DS

VIA VIAG1_E_DS
  LAYER MET5 ;
    RECT -0.200 -0.260 0.320 0.260 ;
  LAYER CUTG1 ;
    RECT -0.140 -0.200 0.260 0.200 ;
  LAYER METG1 ;
    RECT -0.140 -0.200 0.260 0.200 ;
END VIAG1_E_DS

VIA VIAG1_W_DS
  LAYER MET5 ;
    RECT -0.320 -0.260 0.200 0.260 ;
  LAYER CUTG1 ;
    RECT -0.260 -0.200 0.140 0.200 ;
  LAYER METG1 ;
    RECT -0.260 -0.200 0.140 0.200 ;
END VIAG1_W_DS

# MULTI-VIA
VIA VIAG1_2N_DS
  LAYER MET5 ;
    RECT -0.260 -0.260 0.260 1.060 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
    RECT -0.200  0.600 0.200 1.000 ;
  LAYER METG1 ;
    RECT -0.200 -0.200 0.200 1.000 ;
END VIAG1_2N_DS

VIA VIAG1_2S_DS
  LAYER MET5 ;
    RECT -0.260 -1.060 0.260  0.260 ;
  LAYER CUTG1 ;
    RECT -0.200 -1.000 0.200 -0.600 ;
    RECT -0.200 -0.200 0.200  0.200 ;
  LAYER METG1 ;
    RECT -0.200 -1.000 0.200  0.200 ;
END VIAG1_2S_DS

VIA VIAG1_2V_DS
  LAYER MET5 ;
    RECT -0.260 -0.660 0.260  0.660 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.600 0.200 -0.200 ;
    RECT -0.200  0.200 0.200  0.600 ;
  LAYER METG1 ;
    RECT -0.200 -0.600 0.200  0.600 ;
END VIAG1_2V_DS

VIA VIAG1_2E_DS
  LAYER MET5 ;
    RECT -0.260 -0.260 1.060  0.260 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200  0.200 ;
    RECT  0.600 -0.200 1.000  0.200 ;
  LAYER METG1 ;
    RECT -0.200 -0.200 1.000  0.200 ;
END VIAG1_2E_DS

VIA VIAG1_2W_DS
  LAYER MET5 ;
    RECT -1.060 -0.260  0.260 0.260 ;
  LAYER CUTG1 ;
    RECT -1.000 -0.200 -0.600 0.200 ;
    RECT -0.200 -0.200  0.200 0.200 ;
  LAYER METG1 ;
    RECT -1.000 -0.200  0.200 0.200 ;
END VIAG1_2W_DS

VIA VIAG1_2H_DS
  LAYER MET5 ;
    RECT -0.660 -0.260  0.660 0.260 ;
  LAYER CUTG1 ;
    RECT -0.600 -0.200 -0.200 0.200 ;
    RECT  0.200 -0.200  0.600 0.200 ;
  LAYER METG1 ;
    RECT -0.600 -0.200  0.600 0.200 ;
END VIAG1_2H_DS

# SINGLE/STACK-VIA
VIA VIATOP_DS
  LAYER METG1 ;
    RECT -0.350 -0.350 0.350 0.350 ;
  LAYER CUTTOP ;
    RECT -0.250 -0.250 0.250 0.250 ;
  LAYER METTOP ;
    RECT -0.500 -0.500 0.500 0.500 ;
END VIATOP_DS

# MULTI-VIA
VIA VIATOP_2N_DS
  LAYER METG1 ;
    RECT -0.350 -0.350 0.350 1.950 ;
  LAYER CUTTOP ;
    RECT -0.250 -0.250 0.250 0.250 ;
    RECT -0.250  1.350 0.250 1.850 ;
  LAYER METTOP ;
    RECT -0.500 -0.500 0.500 2.100 ;
END VIATOP_2N_DS

VIA VIATOP_2S_DS
  LAYER METG1 ;
    RECT -0.350 -1.950 0.350  0.350 ;
  LAYER CUTTOP ;
    RECT -0.250 -1.850 0.250 -1.350 ;
    RECT -0.250 -0.250 0.250  0.250 ;
  LAYER METTOP ;
    RECT -0.500 -2.100 0.500  0.500 ;
END VIATOP_2S_DS

VIA VIATOP_2V_DS
  LAYER METG1 ;
    RECT -0.350 -1.150 0.350  1.150 ;
  LAYER CUTTOP ;
    RECT -0.250 -1.050 0.250 -0.550 ;
    RECT -0.250  0.550 0.250  1.050 ;
  LAYER METTOP ;
    RECT -0.500 -1.300 0.500  1.300 ;
END VIATOP_2V_DS

VIA VIATOP_2E_DS
  LAYER METG1 ;
    RECT -0.350 -0.350 1.950 0.350 ;
  LAYER CUTTOP ;
    RECT -0.250 -0.250 0.250 0.250 ;
    RECT  1.350 -0.250 1.850 0.250 ;
  LAYER METTOP ;
    RECT -0.500 -0.500 2.100 0.500 ;
END VIATOP_2E_DS

VIA VIATOP_2W_DS
  LAYER METG1 ;
    RECT -1.950 -0.350  0.350 0.350 ;
  LAYER CUTTOP ;
    RECT -1.850 -0.250 -1.350 0.250 ;
    RECT -0.250 -0.250  0.250 0.250 ;
  LAYER METTOP ;
    RECT -2.100 -0.500  0.500 0.500 ;
END VIATOP_2W_DS

VIA VIATOP_2H_DS
  LAYER METG1 ;
    RECT -1.150 -0.350  1.150 0.350 ;
  LAYER CUTTOP ;
    RECT -1.050 -0.250 -0.550 0.250 ;
    RECT  0.550 -0.250  1.050 0.250 ;
  LAYER METTOP ;
    RECT -1.300 -0.500  1.300 0.500 ;
END VIATOP_2H_DS

END DOUBLESPACE

NONDEFAULTRULE DOUBLECUT
LAYER MET1
  WIDTH 0.100 ;
  SPACING 0.100 ;
END MET1

LAYER MET2
  WIDTH 0.100 ;
  SPACING 0.100 ;
END MET2

LAYER MET3
  WIDTH 0.100 ;
  SPACING 0.100 ;
END MET3

LAYER MET4
  WIDTH 0.100 ;
  SPACING 0.100 ;
END MET4

LAYER MET5
  WIDTH 0.100 ;
  SPACING 0.100 ;
END MET5

LAYER METG1
  WIDTH 0.400 ;
  SPACING 0.400 ;
END METG1

LAYER METTOP
  WIDTH 0.800 ;
  SPACING 0.800 ;
END METTOP

# MULTI-VIA
VIA VIA1_2N_MVIA
  LAYER MET1 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA1_2N_MVIA

VIA VIA1_2NV_MVIA
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA1_2NV_MVIA

VIA VIA1_2NR_MVIA
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA1_2NR_MVIA

VIA VIA1_2S_MVIA
  LAYER MET1 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA1_2S_MVIA

VIA VIA1_2SV_MVIA
  LAYER MET1 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA1_2SV_MVIA

VIA VIA1_2SR_MVIA
  LAYER MET1 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA1_2SR_MVIA

VIA VIA1_2V_MVIA
  LAYER MET1 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA1_2V_MVIA

VIA VIA1_2CV_MVIA
  LAYER MET1 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA1_2CV_MVIA

VIA VIA1_2VR_MVIA
  LAYER MET1 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA1_2VR_MVIA

VIA VIA1_2E_MVIA
  LAYER MET1 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA1_2E_MVIA

VIA VIA1_2EH_MVIA
  LAYER MET1 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA1_2EH_MVIA

VIA VIA1_2ER_MVIA
  LAYER MET1 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA1_2ER_MVIA

VIA VIA1_2W_MVIA
  LAYER MET1 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA1_2W_MVIA

VIA VIA1_2WH_MVIA
  LAYER MET1 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA1_2WH_MVIA

VIA VIA1_2WR_MVIA
  LAYER MET1 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA1_2WR_MVIA

VIA VIA1_2H_MVIA
  LAYER MET1 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA1_2H_MVIA

VIA VIA1_2CH_MVIA
  LAYER MET1 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA1_2CH_MVIA

VIA VIA1_2HR_MVIA
  LAYER MET1 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA1_2HR_MVIA

VIA VIA1_3H_MVIA
  LAYER MET1 ;
    RECT -0.290 -0.050  0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.250 -0.090  0.250 0.090 ;
END VIA1_3H_MVIA

VIA VIA1_3V_MVIA
  LAYER MET1 ;
    RECT -0.090 -0.250 0.090  0.250 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.290 ;
END VIA1_3V_MVIA

VIA VIA1_4H_MVIA
  LAYER MET1 ;
    RECT -0.390 -0.050  0.390 0.050 ;
  LAYER CUT12 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET2 ;
    RECT -0.350 -0.090  0.350 0.090 ;
END VIA1_4H_MVIA

VIA VIA1_4V_MVIA
  LAYER MET1 ;
    RECT -0.090 -0.350 0.090  0.350 ;
  LAYER CUT12 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET2 ;
    RECT -0.050 -0.390 0.050  0.390 ;
END VIA1_4V_MVIA

# MULTI-VIA
VIA VIA2_2N_MVIA
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA2_2N_MVIA

VIA VIA2_2NV_MVIA
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA2_2NV_MVIA

VIA VIA2_2NR_MVIA
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA2_2NR_MVIA

VIA VIA2_2S_MVIA
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA2_2S_MVIA

VIA VIA2_2SV_MVIA
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA2_2SV_MVIA

VIA VIA2_2SR_MVIA
  LAYER MET2 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA2_2SR_MVIA

VIA VIA2_2V_MVIA
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA2_2V_MVIA

VIA VIA2_2CV_MVIA
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA2_2CV_MVIA

VIA VIA2_2VR_MVIA
  LAYER MET2 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA2_2VR_MVIA

VIA VIA2_2E_MVIA
  LAYER MET2 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA2_2E_MVIA

VIA VIA2_2EH_MVIA
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA2_2EH_MVIA

VIA VIA2_2ER_MVIA
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA2_2ER_MVIA

VIA VIA2_2W_MVIA
  LAYER MET2 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA2_2W_MVIA

VIA VIA2_2WH_MVIA
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA2_2WH_MVIA

VIA VIA2_2WR_MVIA
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA2_2WR_MVIA

VIA VIA2_2H_MVIA
  LAYER MET2 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA2_2H_MVIA

VIA VIA2_2CH_MVIA
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA2_2CH_MVIA

VIA VIA2_2HR_MVIA
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA2_2HR_MVIA

VIA VIA2_3H_MVIA
  LAYER MET2 ;
    RECT -0.250 -0.090  0.250 0.090 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.290 0.050 ;
END VIA2_3H_MVIA

VIA VIA2_3V_MVIA
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.250 ;
END VIA2_3V_MVIA

VIA VIA2_4H_MVIA
  LAYER MET2 ;
    RECT -0.350 -0.090  0.350 0.090 ;
  LAYER CUT23 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET3 ;
    RECT -0.390 -0.050  0.390 0.050 ;
END VIA2_4H_MVIA

VIA VIA2_4V_MVIA
  LAYER MET2 ;
    RECT -0.050 -0.390 0.050  0.390 ;
  LAYER CUT23 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET3 ;
    RECT -0.090 -0.350 0.090  0.350 ;
END VIA2_4V_MVIA

# MULTI-VIA
VIA VIA3_2N_MVIA
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA3_2N_MVIA

VIA VIA3_2NV_MVIA
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA3_2NV_MVIA

VIA VIA3_2NR_MVIA
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA3_2NR_MVIA

VIA VIA3_2S_MVIA
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA3_2S_MVIA

VIA VIA3_2SV_MVIA
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA3_2SV_MVIA

VIA VIA3_2SR_MVIA
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA3_2SR_MVIA

VIA VIA3_2V_MVIA
  LAYER MET3 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT34 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA3_2V_MVIA

VIA VIA3_2CV_MVIA
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT34 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA3_2CV_MVIA

VIA VIA3_2VR_MVIA
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT34 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET4 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA3_2VR_MVIA

VIA VIA3_2E_MVIA
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA3_2E_MVIA

VIA VIA3_2EH_MVIA
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA3_2EH_MVIA

VIA VIA3_2ER_MVIA
  LAYER MET3 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA3_2ER_MVIA

VIA VIA3_2W_MVIA
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA3_2W_MVIA

VIA VIA3_2WH_MVIA
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA3_2WH_MVIA

VIA VIA3_2WR_MVIA
  LAYER MET3 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA3_2WR_MVIA

VIA VIA3_2H_MVIA
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT34 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET4 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA3_2H_MVIA

VIA VIA3_2CH_MVIA
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT34 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET4 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA3_2CH_MVIA

VIA VIA3_2HR_MVIA
  LAYER MET3 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT34 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET4 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA3_2HR_MVIA

VIA VIA3_3H_MVIA
  LAYER MET3 ;
    RECT -0.290 -0.050  0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.250 -0.090  0.250 0.090 ;
END VIA3_3H_MVIA

VIA VIA3_3V_MVIA
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.250 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.290 ;
END VIA3_3V_MVIA

VIA VIA3_4H_MVIA
  LAYER MET3 ;
    RECT -0.390 -0.050  0.390 0.050 ;
  LAYER CUT34 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET4 ;
    RECT -0.350 -0.090  0.350 0.090 ;
END VIA3_4H_MVIA

VIA VIA3_4V_MVIA
  LAYER MET3 ;
    RECT -0.090 -0.350 0.090  0.350 ;
  LAYER CUT34 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET4 ;
    RECT -0.050 -0.390 0.050  0.390 ;
END VIA3_4V_MVIA

# MULTI-VIA
VIA VIA4_2N_MVIA
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA4_2N_MVIA

VIA VIA4_2NV_MVIA
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA4_2NV_MVIA

VIA VIA4_2NR_MVIA
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA4_2NR_MVIA

VIA VIA4_2S_MVIA
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA4_2S_MVIA

VIA VIA4_2SV_MVIA
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA4_2SV_MVIA

VIA VIA4_2SR_MVIA
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA4_2SR_MVIA

VIA VIA4_2V_MVIA
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT45 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET5 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA4_2V_MVIA

VIA VIA4_2CV_MVIA
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT45 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET5 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA4_2CV_MVIA

VIA VIA4_2VR_MVIA
  LAYER MET4 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT45 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET5 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA4_2VR_MVIA

VIA VIA4_2E_MVIA
  LAYER MET4 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA4_2E_MVIA

VIA VIA4_2EH_MVIA
  LAYER MET4 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA4_2EH_MVIA

VIA VIA4_2ER_MVIA
  LAYER MET4 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA4_2ER_MVIA

VIA VIA4_2W_MVIA
  LAYER MET4 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA4_2W_MVIA

VIA VIA4_2WH_MVIA
  LAYER MET4 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA4_2WH_MVIA

VIA VIA4_2WR_MVIA
  LAYER MET4 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA4_2WR_MVIA

VIA VIA4_2H_MVIA
  LAYER MET4 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT45 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET5 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA4_2H_MVIA

VIA VIA4_2CH_MVIA
  LAYER MET4 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT45 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET5 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA4_2CH_MVIA

VIA VIA4_2HR_MVIA
  LAYER MET4 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT45 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET5 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA4_2HR_MVIA

VIA VIA4_3H_MVIA
  LAYER MET4 ;
    RECT -0.250 -0.090  0.250 0.090 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.290 -0.050  0.290 0.050 ;
END VIA4_3H_MVIA

VIA VIA4_3V_MVIA
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.290 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET5 ;
    RECT -0.090 -0.250 0.090  0.250 ;
END VIA4_3V_MVIA

VIA VIA4_4H_MVIA
  LAYER MET4 ;
    RECT -0.350 -0.090  0.350 0.090 ;
  LAYER CUT45 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET5 ;
    RECT -0.390 -0.050  0.390 0.050 ;
END VIA4_4H_MVIA

VIA VIA4_4V_MVIA
  LAYER MET4 ;
    RECT -0.050 -0.390 0.050  0.390 ;
  LAYER CUT45 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET5 ;
    RECT -0.090 -0.350 0.090  0.350 ;
END VIA4_4V_MVIA

# MULTI-VIA
VIA VIAG1_2N_MVIA
  LAYER MET5 ;
    RECT -0.260 -0.260 0.260 1.060 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
    RECT -0.200  0.600 0.200 1.000 ;
  LAYER METG1 ;
    RECT -0.200 -0.200 0.200 1.000 ;
END VIAG1_2N_MVIA

VIA VIAG1_2S_MVIA
  LAYER MET5 ;
    RECT -0.260 -1.060 0.260  0.260 ;
  LAYER CUTG1 ;
    RECT -0.200 -1.000 0.200 -0.600 ;
    RECT -0.200 -0.200 0.200  0.200 ;
  LAYER METG1 ;
    RECT -0.200 -1.000 0.200  0.200 ;
END VIAG1_2S_MVIA

VIA VIAG1_2V_MVIA
  LAYER MET5 ;
    RECT -0.260 -0.660 0.260  0.660 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.600 0.200 -0.200 ;
    RECT -0.200  0.200 0.200  0.600 ;
  LAYER METG1 ;
    RECT -0.200 -0.600 0.200  0.600 ;
END VIAG1_2V_MVIA

VIA VIAG1_2E_MVIA
  LAYER MET5 ;
    RECT -0.260 -0.260 1.060  0.260 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200  0.200 ;
    RECT  0.600 -0.200 1.000  0.200 ;
  LAYER METG1 ;
    RECT -0.200 -0.200 1.000  0.200 ;
END VIAG1_2E_MVIA

VIA VIAG1_2W_MVIA
  LAYER MET5 ;
    RECT -1.060 -0.260  0.260 0.260 ;
  LAYER CUTG1 ;
    RECT -1.000 -0.200 -0.600 0.200 ;
    RECT -0.200 -0.200  0.200 0.200 ;
  LAYER METG1 ;
    RECT -1.000 -0.200  0.200 0.200 ;
END VIAG1_2W_MVIA

VIA VIAG1_2H_MVIA
  LAYER MET5 ;
    RECT -0.660 -0.260  0.660 0.260 ;
  LAYER CUTG1 ;
    RECT -0.600 -0.200 -0.200 0.200 ;
    RECT  0.200 -0.200  0.600 0.200 ;
  LAYER METG1 ;
    RECT -0.600 -0.200  0.600 0.200 ;
END VIAG1_2H_MVIA

# MULTI-VIA
VIA VIATOP_2N_MVIA
  LAYER METG1 ;
    RECT -0.350 -0.350 0.350 1.950 ;
  LAYER CUTTOP ;
    RECT -0.250 -0.250 0.250 0.250 ;
    RECT -0.250  1.350 0.250 1.850 ;
  LAYER METTOP ;
    RECT -0.500 -0.500 0.500 2.100 ;
END VIATOP_2N_MVIA

VIA VIATOP_2S_MVIA
  LAYER METG1 ;
    RECT -0.350 -1.950 0.350  0.350 ;
  LAYER CUTTOP ;
    RECT -0.250 -1.850 0.250 -1.350 ;
    RECT -0.250 -0.250 0.250  0.250 ;
  LAYER METTOP ;
    RECT -0.500 -2.100 0.500  0.500 ;
END VIATOP_2S_MVIA

VIA VIATOP_2V_MVIA
  LAYER METG1 ;
    RECT -0.350 -1.150 0.350  1.150 ;
  LAYER CUTTOP ;
    RECT -0.250 -1.050 0.250 -0.550 ;
    RECT -0.250  0.550 0.250  1.050 ;
  LAYER METTOP ;
    RECT -0.500 -1.300 0.500  1.300 ;
END VIATOP_2V_MVIA

VIA VIATOP_2E_MVIA
  LAYER METG1 ;
    RECT -0.350 -0.350 1.950 0.350 ;
  LAYER CUTTOP ;
    RECT -0.250 -0.250 0.250 0.250 ;
    RECT  1.350 -0.250 1.850 0.250 ;
  LAYER METTOP ;
    RECT -0.500 -0.500 2.100 0.500 ;
END VIATOP_2E_MVIA

VIA VIATOP_2W_MVIA
  LAYER METG1 ;
    RECT -1.950 -0.350  0.350 0.350 ;
  LAYER CUTTOP ;
    RECT -1.850 -0.250 -1.350 0.250 ;
    RECT -0.250 -0.250  0.250 0.250 ;
  LAYER METTOP ;
    RECT -2.100 -0.500  0.500 0.500 ;
END VIATOP_2W_MVIA

VIA VIATOP_2H_MVIA
  LAYER METG1 ;
    RECT -1.150 -0.350  1.150 0.350 ;
  LAYER CUTTOP ;
    RECT -1.050 -0.250 -0.550 0.250 ;
    RECT  0.550 -0.250  1.050 0.250 ;
  LAYER METTOP ;
    RECT -1.300 -0.500  1.300 0.500 ;
END VIATOP_2H_MVIA

END DOUBLECUT

NONDEFAULTRULE DOUBLECUT_DS
LAYER MET1
  WIDTH 0.100 ;
  SPACING 0.200 ;
END MET1

LAYER MET2
  WIDTH 0.100 ;
  SPACING 0.200 ;
END MET2

LAYER MET3
  WIDTH 0.100 ;
  SPACING 0.200 ;
END MET3

LAYER MET4
  WIDTH 0.100 ;
  SPACING 0.200 ;
END MET4

LAYER MET5
  WIDTH 0.100 ;
  SPACING 0.200 ;
END MET5

LAYER METG1
  WIDTH 0.400 ;
  SPACING 0.800 ;
END METG1

LAYER METTOP
  WIDTH 0.800 ;
  SPACING 1.600 ;
END METTOP

# MULTI-VIA
VIA VIA1_2N_DSMVIA
  LAYER MET1 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA1_2N_DSMVIA

VIA VIA1_2NV_DSMVIA
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA1_2NV_DSMVIA

VIA VIA1_2NR_DSMVIA
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA1_2NR_DSMVIA

VIA VIA1_2S_DSMVIA
  LAYER MET1 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA1_2S_DSMVIA

VIA VIA1_2SV_DSMVIA
  LAYER MET1 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA1_2SV_DSMVIA

VIA VIA1_2SR_DSMVIA
  LAYER MET1 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA1_2SR_DSMVIA

VIA VIA1_2V_DSMVIA
  LAYER MET1 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA1_2V_DSMVIA

VIA VIA1_2CV_DSMVIA
  LAYER MET1 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA1_2CV_DSMVIA

VIA VIA1_2VR_DSMVIA
  LAYER MET1 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA1_2VR_DSMVIA

VIA VIA1_2E_DSMVIA
  LAYER MET1 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA1_2E_DSMVIA

VIA VIA1_2EH_DSMVIA
  LAYER MET1 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA1_2EH_DSMVIA

VIA VIA1_2ER_DSMVIA
  LAYER MET1 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA1_2ER_DSMVIA

VIA VIA1_2W_DSMVIA
  LAYER MET1 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA1_2W_DSMVIA

VIA VIA1_2WH_DSMVIA
  LAYER MET1 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA1_2WH_DSMVIA

VIA VIA1_2WR_DSMVIA
  LAYER MET1 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA1_2WR_DSMVIA

VIA VIA1_2H_DSMVIA
  LAYER MET1 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA1_2H_DSMVIA

VIA VIA1_2CH_DSMVIA
  LAYER MET1 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA1_2CH_DSMVIA

VIA VIA1_2HR_DSMVIA
  LAYER MET1 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA1_2HR_DSMVIA

VIA VIA1_3H_DSMVIA
  LAYER MET1 ;
    RECT -0.290 -0.050  0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.250 -0.090  0.250 0.090 ;
END VIA1_3H_DSMVIA

VIA VIA1_3V_DSMVIA
  LAYER MET1 ;
    RECT -0.090 -0.250 0.090  0.250 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.290 ;
END VIA1_3V_DSMVIA

VIA VIA1_4H_DSMVIA
  LAYER MET1 ;
    RECT -0.390 -0.050  0.390 0.050 ;
  LAYER CUT12 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET2 ;
    RECT -0.350 -0.090  0.350 0.090 ;
END VIA1_4H_DSMVIA

VIA VIA1_4V_DSMVIA
  LAYER MET1 ;
    RECT -0.090 -0.350 0.090  0.350 ;
  LAYER CUT12 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET2 ;
    RECT -0.050 -0.390 0.050  0.390 ;
END VIA1_4V_DSMVIA

# MULTI-VIA
VIA VIA2_2N_DSMVIA
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA2_2N_DSMVIA

VIA VIA2_2NV_DSMVIA
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA2_2NV_DSMVIA

VIA VIA2_2NR_DSMVIA
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA2_2NR_DSMVIA

VIA VIA2_2S_DSMVIA
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA2_2S_DSMVIA

VIA VIA2_2SV_DSMVIA
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA2_2SV_DSMVIA

VIA VIA2_2SR_DSMVIA
  LAYER MET2 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA2_2SR_DSMVIA

VIA VIA2_2V_DSMVIA
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA2_2V_DSMVIA

VIA VIA2_2CV_DSMVIA
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA2_2CV_DSMVIA

VIA VIA2_2VR_DSMVIA
  LAYER MET2 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA2_2VR_DSMVIA

VIA VIA2_2E_DSMVIA
  LAYER MET2 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA2_2E_DSMVIA

VIA VIA2_2EH_DSMVIA
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA2_2EH_DSMVIA

VIA VIA2_2ER_DSMVIA
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA2_2ER_DSMVIA

VIA VIA2_2W_DSMVIA
  LAYER MET2 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA2_2W_DSMVIA

VIA VIA2_2WH_DSMVIA
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA2_2WH_DSMVIA

VIA VIA2_2WR_DSMVIA
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA2_2WR_DSMVIA

VIA VIA2_2H_DSMVIA
  LAYER MET2 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA2_2H_DSMVIA

VIA VIA2_2CH_DSMVIA
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA2_2CH_DSMVIA

VIA VIA2_2HR_DSMVIA
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA2_2HR_DSMVIA

VIA VIA2_3H_DSMVIA
  LAYER MET2 ;
    RECT -0.250 -0.090  0.250 0.090 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.290 0.050 ;
END VIA2_3H_DSMVIA

VIA VIA2_3V_DSMVIA
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.250 ;
END VIA2_3V_DSMVIA

VIA VIA2_4H_DSMVIA
  LAYER MET2 ;
    RECT -0.350 -0.090  0.350 0.090 ;
  LAYER CUT23 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET3 ;
    RECT -0.390 -0.050  0.390 0.050 ;
END VIA2_4H_DSMVIA

VIA VIA2_4V_DSMVIA
  LAYER MET2 ;
    RECT -0.050 -0.390 0.050  0.390 ;
  LAYER CUT23 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET3 ;
    RECT -0.090 -0.350 0.090  0.350 ;
END VIA2_4V_DSMVIA

# MULTI-VIA
VIA VIA3_2N_DSMVIA
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA3_2N_DSMVIA

VIA VIA3_2NV_DSMVIA
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA3_2NV_DSMVIA

VIA VIA3_2NR_DSMVIA
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA3_2NR_DSMVIA

VIA VIA3_2S_DSMVIA
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA3_2S_DSMVIA

VIA VIA3_2SV_DSMVIA
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA3_2SV_DSMVIA

VIA VIA3_2SR_DSMVIA
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA3_2SR_DSMVIA

VIA VIA3_2V_DSMVIA
  LAYER MET3 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT34 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA3_2V_DSMVIA

VIA VIA3_2CV_DSMVIA
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT34 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA3_2CV_DSMVIA

VIA VIA3_2VR_DSMVIA
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT34 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET4 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA3_2VR_DSMVIA

VIA VIA3_2E_DSMVIA
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA3_2E_DSMVIA

VIA VIA3_2EH_DSMVIA
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA3_2EH_DSMVIA

VIA VIA3_2ER_DSMVIA
  LAYER MET3 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA3_2ER_DSMVIA

VIA VIA3_2W_DSMVIA
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA3_2W_DSMVIA

VIA VIA3_2WH_DSMVIA
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA3_2WH_DSMVIA

VIA VIA3_2WR_DSMVIA
  LAYER MET3 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA3_2WR_DSMVIA

VIA VIA3_2H_DSMVIA
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT34 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET4 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA3_2H_DSMVIA

VIA VIA3_2CH_DSMVIA
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT34 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET4 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA3_2CH_DSMVIA

VIA VIA3_2HR_DSMVIA
  LAYER MET3 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT34 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET4 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA3_2HR_DSMVIA

VIA VIA3_3H_DSMVIA
  LAYER MET3 ;
    RECT -0.290 -0.050  0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.250 -0.090  0.250 0.090 ;
END VIA3_3H_DSMVIA

VIA VIA3_3V_DSMVIA
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.250 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.290 ;
END VIA3_3V_DSMVIA

VIA VIA3_4H_DSMVIA
  LAYER MET3 ;
    RECT -0.390 -0.050  0.390 0.050 ;
  LAYER CUT34 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET4 ;
    RECT -0.350 -0.090  0.350 0.090 ;
END VIA3_4H_DSMVIA

VIA VIA3_4V_DSMVIA
  LAYER MET3 ;
    RECT -0.090 -0.350 0.090  0.350 ;
  LAYER CUT34 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET4 ;
    RECT -0.050 -0.390 0.050  0.390 ;
END VIA3_4V_DSMVIA

# MULTI-VIA
VIA VIA4_2N_DSMVIA
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA4_2N_DSMVIA

VIA VIA4_2NV_DSMVIA
  LAYER MET4 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA4_2NV_DSMVIA

VIA VIA4_2NR_DSMVIA
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA4_2NR_DSMVIA

VIA VIA4_2S_DSMVIA
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA4_2S_DSMVIA

VIA VIA4_2SV_DSMVIA
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA4_2SV_DSMVIA

VIA VIA4_2SR_DSMVIA
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA4_2SR_DSMVIA

VIA VIA4_2V_DSMVIA
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT45 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET5 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA4_2V_DSMVIA

VIA VIA4_2CV_DSMVIA
  LAYER MET4 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT45 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET5 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA4_2CV_DSMVIA

VIA VIA4_2VR_DSMVIA
  LAYER MET4 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT45 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET5 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA4_2VR_DSMVIA

VIA VIA4_2E_DSMVIA
  LAYER MET4 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA4_2E_DSMVIA

VIA VIA4_2EH_DSMVIA
  LAYER MET4 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA4_2EH_DSMVIA

VIA VIA4_2ER_DSMVIA
  LAYER MET4 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA4_2ER_DSMVIA

VIA VIA4_2W_DSMVIA
  LAYER MET4 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA4_2W_DSMVIA

VIA VIA4_2WH_DSMVIA
  LAYER MET4 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA4_2WH_DSMVIA

VIA VIA4_2WR_DSMVIA
  LAYER MET4 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA4_2WR_DSMVIA

VIA VIA4_2H_DSMVIA
  LAYER MET4 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT45 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET5 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA4_2H_DSMVIA

VIA VIA4_2CH_DSMVIA
  LAYER MET4 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT45 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET5 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA4_2CH_DSMVIA

VIA VIA4_2HR_DSMVIA
  LAYER MET4 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT45 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET5 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA4_2HR_DSMVIA

VIA VIA4_3H_DSMVIA
  LAYER MET4 ;
    RECT -0.250 -0.090  0.250 0.090 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.290 -0.050  0.290 0.050 ;
END VIA4_3H_DSMVIA

VIA VIA4_3V_DSMVIA
  LAYER MET4 ;
    RECT -0.050 -0.290 0.050  0.290 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET5 ;
    RECT -0.090 -0.250 0.090  0.250 ;
END VIA4_3V_DSMVIA

VIA VIA4_4H_DSMVIA
  LAYER MET4 ;
    RECT -0.350 -0.090  0.350 0.090 ;
  LAYER CUT45 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET5 ;
    RECT -0.390 -0.050  0.390 0.050 ;
END VIA4_4H_DSMVIA

VIA VIA4_4V_DSMVIA
  LAYER MET4 ;
    RECT -0.050 -0.390 0.050  0.390 ;
  LAYER CUT45 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET5 ;
    RECT -0.090 -0.350 0.090  0.350 ;
END VIA4_4V_DSMVIA

# MULTI-VIA
VIA VIAG1_2N_DSMVIA
  LAYER MET5 ;
    RECT -0.260 -0.260 0.260 1.060 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
    RECT -0.200  0.600 0.200 1.000 ;
  LAYER METG1 ;
    RECT -0.200 -0.200 0.200 1.000 ;
END VIAG1_2N_DSMVIA

VIA VIAG1_2S_DSMVIA
  LAYER MET5 ;
    RECT -0.260 -1.060 0.260  0.260 ;
  LAYER CUTG1 ;
    RECT -0.200 -1.000 0.200 -0.600 ;
    RECT -0.200 -0.200 0.200  0.200 ;
  LAYER METG1 ;
    RECT -0.200 -1.000 0.200  0.200 ;
END VIAG1_2S_DSMVIA

VIA VIAG1_2V_DSMVIA
  LAYER MET5 ;
    RECT -0.260 -0.660 0.260  0.660 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.600 0.200 -0.200 ;
    RECT -0.200  0.200 0.200  0.600 ;
  LAYER METG1 ;
    RECT -0.200 -0.600 0.200  0.600 ;
END VIAG1_2V_DSMVIA

VIA VIAG1_2E_DSMVIA
  LAYER MET5 ;
    RECT -0.260 -0.260 1.060  0.260 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200  0.200 ;
    RECT  0.600 -0.200 1.000  0.200 ;
  LAYER METG1 ;
    RECT -0.200 -0.200 1.000  0.200 ;
END VIAG1_2E_DSMVIA

VIA VIAG1_2W_DSMVIA
  LAYER MET5 ;
    RECT -1.060 -0.260  0.260 0.260 ;
  LAYER CUTG1 ;
    RECT -1.000 -0.200 -0.600 0.200 ;
    RECT -0.200 -0.200  0.200 0.200 ;
  LAYER METG1 ;
    RECT -1.000 -0.200  0.200 0.200 ;
END VIAG1_2W_DSMVIA

VIA VIAG1_2H_DSMVIA
  LAYER MET5 ;
    RECT -0.660 -0.260  0.660 0.260 ;
  LAYER CUTG1 ;
    RECT -0.600 -0.200 -0.200 0.200 ;
    RECT  0.200 -0.200  0.600 0.200 ;
  LAYER METG1 ;
    RECT -0.600 -0.200  0.600 0.200 ;
END VIAG1_2H_DSMVIA

# MULTI-VIA
VIA VIATOP_2N_DSMVIA
  LAYER METG1 ;
    RECT -0.350 -0.350 0.350 1.950 ;
  LAYER CUTTOP ;
    RECT -0.250 -0.250 0.250 0.250 ;
    RECT -0.250  1.350 0.250 1.850 ;
  LAYER METTOP ;
    RECT -0.500 -0.500 0.500 2.100 ;
END VIATOP_2N_DSMVIA

VIA VIATOP_2S_DSMVIA
  LAYER METG1 ;
    RECT -0.350 -1.950 0.350  0.350 ;
  LAYER CUTTOP ;
    RECT -0.250 -1.850 0.250 -1.350 ;
    RECT -0.250 -0.250 0.250  0.250 ;
  LAYER METTOP ;
    RECT -0.500 -2.100 0.500  0.500 ;
END VIATOP_2S_DSMVIA

VIA VIATOP_2V_DSMVIA
  LAYER METG1 ;
    RECT -0.350 -1.150 0.350  1.150 ;
  LAYER CUTTOP ;
    RECT -0.250 -1.050 0.250 -0.550 ;
    RECT -0.250  0.550 0.250  1.050 ;
  LAYER METTOP ;
    RECT -0.500 -1.300 0.500  1.300 ;
END VIATOP_2V_DSMVIA

VIA VIATOP_2E_DSMVIA
  LAYER METG1 ;
    RECT -0.350 -0.350 1.950 0.350 ;
  LAYER CUTTOP ;
    RECT -0.250 -0.250 0.250 0.250 ;
    RECT  1.350 -0.250 1.850 0.250 ;
  LAYER METTOP ;
    RECT -0.500 -0.500 2.100 0.500 ;
END VIATOP_2E_DSMVIA

VIA VIATOP_2W_DSMVIA
  LAYER METG1 ;
    RECT -1.950 -0.350  0.350 0.350 ;
  LAYER CUTTOP ;
    RECT -1.850 -0.250 -1.350 0.250 ;
    RECT -0.250 -0.250  0.250 0.250 ;
  LAYER METTOP ;
    RECT -2.100 -0.500  0.500 0.500 ;
END VIATOP_2W_DSMVIA

VIA VIATOP_2H_DSMVIA
  LAYER METG1 ;
    RECT -1.150 -0.350  1.150 0.350 ;
  LAYER CUTTOP ;
    RECT -1.050 -0.250 -0.550 0.250 ;
    RECT  0.550 -0.250  1.050 0.250 ;
  LAYER METTOP ;
    RECT -1.300 -0.500  1.300 0.500 ;
END VIATOP_2H_DSMVIA

END DOUBLECUT_DS

NONDEFAULTRULE WIDEWIRE
LAYER MET1
  WIDTH 0.100 ;
  SPACING 0.100 ;
END MET1

LAYER MET2
  WIDTH 0.100 ;
  SPACING 0.100 ;
END MET2

LAYER MET3
  WIDTH 0.100 ;
  SPACING 0.100 ;
END MET3

LAYER MET4
  WIDTH 0.180 ;
  SPACING 0.120 ;
END MET4

LAYER MET5
  WIDTH 0.180 ;
  SPACING 0.120 ;
END MET5

LAYER METG1
  WIDTH 0.400 ;
  SPACING 0.400 ;
END METG1

LAYER METTOP
  WIDTH 0.800 ;
  SPACING 0.800 ;
END METTOP

# SINGLE-VIA
VIA VIA1_HV_WW
  LAYER MET1 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA1_HV_WW

VIA VIA1_HH_WW
  LAYER MET1 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA1_HH_WW

VIA VIA1_VH_WW
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA1_VH_WW

VIA VIA1_VV_WW
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA1_VV_WW

# MULTI-VIA
VIA VIA1_2N_WW
  LAYER MET1 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA1_2N_WW

VIA VIA1_2NV_WW
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA1_2NV_WW

VIA VIA1_2NR_WW
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA1_2NR_WW

VIA VIA1_2S_WW
  LAYER MET1 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA1_2S_WW

VIA VIA1_2SV_WW
  LAYER MET1 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA1_2SV_WW

VIA VIA1_2SR_WW
  LAYER MET1 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA1_2SR_WW

VIA VIA1_2V_WW
  LAYER MET1 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA1_2V_WW

VIA VIA1_2CV_WW
  LAYER MET1 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA1_2CV_WW

VIA VIA1_2VR_WW
  LAYER MET1 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA1_2VR_WW

VIA VIA1_2E_WW
  LAYER MET1 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA1_2E_WW

VIA VIA1_2EH_WW
  LAYER MET1 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA1_2EH_WW

VIA VIA1_2ER_WW
  LAYER MET1 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA1_2ER_WW

VIA VIA1_2W_WW
  LAYER MET1 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA1_2W_WW

VIA VIA1_2WH_WW
  LAYER MET1 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA1_2WH_WW

VIA VIA1_2WR_WW
  LAYER MET1 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA1_2WR_WW

VIA VIA1_2H_WW
  LAYER MET1 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA1_2H_WW

VIA VIA1_2CH_WW
  LAYER MET1 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA1_2CH_WW

VIA VIA1_2HR_WW
  LAYER MET1 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA1_2HR_WW

VIA VIA1_3H_WW
  LAYER MET1 ;
    RECT -0.290 -0.050  0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.250 -0.090  0.250 0.090 ;
END VIA1_3H_WW

VIA VIA1_3V_WW
  LAYER MET1 ;
    RECT -0.090 -0.250 0.090  0.250 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.290 ;
END VIA1_3V_WW

VIA VIA1_4H_WW
  LAYER MET1 ;
    RECT -0.390 -0.050  0.390 0.050 ;
  LAYER CUT12 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET2 ;
    RECT -0.350 -0.090  0.350 0.090 ;
END VIA1_4H_WW

VIA VIA1_4V_WW
  LAYER MET1 ;
    RECT -0.090 -0.350 0.090  0.350 ;
  LAYER CUT12 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET2 ;
    RECT -0.050 -0.390 0.050  0.390 ;
END VIA1_4V_WW

# SINGLE-VIA
VIA VIA2_VH_WW
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA2_VH_WW

VIA VIA2_VV_WW
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA2_VV_WW

VIA VIA2_HV_WW
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.090 ;
END VIA2_HV_WW

VIA VIA2_HH_WW
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA2_HH_WW

# STACK-VIA
VIA VIA2_NS_WW
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA2_NS_WW

VIA VIA2_SS_WW
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050 0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA2_SS_WW

VIA VIA2_VS_WW
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050 0.190 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
END VIA2_VS_WW

# MULTI-VIA
VIA VIA2_2N_WW
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA2_2N_WW

VIA VIA2_2S_WW
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA2_2S_WW

VIA VIA2_2V_WW
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA2_2V_WW

VIA VIA2_2E_WW
  LAYER MET2 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA2_2E_WW

VIA VIA2_2W_WW
  LAYER MET2 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA2_2W_WW

VIA VIA2_2H_WW
  LAYER MET2 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA2_2H_WW

VIA VIA2_2NR_WW
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA2_2NR_WW

VIA VIA2_2SR_WW
  LAYER MET2 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA2_2SR_WW

VIA VIA2_2VR_WW
  LAYER MET2 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA2_2VR_WW

VIA VIA2_2ER_WW
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA2_2ER_WW

VIA VIA2_2WR_WW
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA2_2WR_WW

VIA VIA2_2HR_WW
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA2_2HR_WW

VIA VIA2_2NV_WW
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA2_2NV_WW

VIA VIA2_2SV_WW
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA2_2SV_WW

VIA VIA2_2CV_WW
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA2_2CV_WW

VIA VIA2_2EH_WW
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA2_2EH_WW

VIA VIA2_2WH_WW
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA2_2WH_WW

VIA VIA2_2CH_WW
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA2_2CH_WW

VIA VIA2_3H_WW
  LAYER MET2 ;
    RECT -0.250 -0.090  0.250 0.090 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.290 0.050 ;
END VIA2_3H_WW

VIA VIA2_3V_WW
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.250 ;
END VIA2_3V_WW

VIA VIA2_4H_WW
  LAYER MET2 ;
    RECT -0.350 -0.090  0.350 0.090 ;
  LAYER CUT23 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET3 ;
    RECT -0.390 -0.050  0.390 0.050 ;
END VIA2_4H_WW

VIA VIA2_4V_WW
  LAYER MET2 ;
    RECT -0.050 -0.390 0.050  0.390 ;
  LAYER CUT23 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET3 ;
    RECT -0.090 -0.350 0.090  0.350 ;
END VIA2_4V_WW

# SINGLE-VIA
VIA VIA3_H_WW
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.090 0.090 0.090 ;
END VIA3_H_WW

VIA VIA3_V_WW
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.090 0.090 0.090 ;
END VIA3_V_WW

# STACK-VIA
VIA VIA3_ES_WW
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.090 0.090 0.090 ;
END VIA3_ES_WW

VIA VIA3_WS_WW
  LAYER MET3 ;
    RECT -0.290 -0.050 0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.090 0.090 0.090 ;
END VIA3_WS_WW

VIA VIA3_HS_WW
  LAYER MET3 ;
    RECT -0.190 -0.050 0.190 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.090 0.090 0.090 ;
END VIA3_HS_WW

# MULTI-VIA
VIA VIA3_2N_WW
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA3_2N_WW

VIA VIA3_2S_WW
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA3_2S_WW

VIA VIA3_2E_WW
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA3_2E_WW

VIA VIA3_2W_WW
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA3_2W_WW

VIA VIA3_2NR_WW
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA3_2NR_WW

VIA VIA3_2SR_WW
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA3_2SR_WW

VIA VIA3_2ER_WW
  LAYER MET3 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA3_2ER_WW

VIA VIA3_2WR_WW
  LAYER MET3 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA3_2WR_WW

VIA VIA3_2CH_WW
  LAYER MET3 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT34 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET4 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA3_2CH_WW

VIA VIA3_2VR_WW
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT34 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET4 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA3_2VR_WW

VIA VIA3_3H_WW
  LAYER MET3 ;
    RECT -0.290 -0.050  0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.250 -0.090  0.250 0.090 ;
END VIA3_3H_WW

VIA VIA3_3V_WW
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.250 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.250 ;
END VIA3_3V_WW

VIA VIA3_4H_WW
  LAYER MET3 ;
    RECT -0.390 -0.050  0.390 0.050 ;
  LAYER CUT34 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET4 ;
    RECT -0.350 -0.090  0.350 0.090 ;
END VIA3_4H_WW

VIA VIA3_4V_WW
  LAYER MET3 ;
    RECT -0.090 -0.350 0.090  0.350 ;
  LAYER CUT34 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET4 ;
    RECT -0.090 -0.350 0.090  0.350 ;
END VIA3_4V_WW

# SINGLE-VIA
VIA VIA4__WW
  LAYER MET4 ;
    RECT -0.090 -0.090 0.090 0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.090 0.090 0.090 ;
END VIA4__WW

# STACK-VIA
VIA VIA4_NS_WW
  LAYER MET4 ;
    RECT -0.090 -0.090 0.090 0.130 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.090 0.090 0.090 ;
END VIA4_NS_WW

VIA VIA4_SS_WW
  LAYER MET4 ;
    RECT -0.090 -0.130 0.090 0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.090 0.090 0.090 ;
END VIA4_SS_WW

VIA VIA4_VS_WW
  LAYER MET4 ;
    RECT -0.090 -0.110 0.090 0.110 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.090 0.090 0.090 ;
END VIA4_VS_WW

# MULTI-VIA
VIA VIA4_2N_WW
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA4_2N_WW

VIA VIA4_2S_WW
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA4_2S_WW

VIA VIA4_2V_WW
  LAYER MET4 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT45 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET5 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA4_2V_WW

VIA VIA4_2E_WW
  LAYER MET4 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA4_2E_WW

VIA VIA4_2W_WW
  LAYER MET4 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA4_2W_WW

VIA VIA4_2H_WW
  LAYER MET4 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT45 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET5 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA4_2H_WW

VIA VIA4_3H_WW
  LAYER MET4 ;
    RECT -0.250 -0.090  0.250 0.090 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.250 -0.090  0.250 0.090 ;
END VIA4_3H_WW

VIA VIA4_3V_WW
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.250 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET5 ;
    RECT -0.090 -0.250 0.090  0.250 ;
END VIA4_3V_WW

VIA VIA4_4H_WW
  LAYER MET4 ;
    RECT -0.350 -0.090  0.350 0.090 ;
  LAYER CUT45 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET5 ;
    RECT -0.350 -0.090  0.350 0.090 ;
END VIA4_4H_WW

VIA VIA4_4V_WW
  LAYER MET4 ;
    RECT -0.090 -0.350 0.090  0.350 ;
  LAYER CUT45 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET5 ;
    RECT -0.090 -0.350 0.090  0.350 ;
END VIA4_4V_WW

# SINGLE/STACK-VIA
VIA VIAG1_WW
  LAYER MET5 ;
    RECT -0.260 -0.260 0.260 0.260 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
  LAYER METG1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
END VIAG1_WW

VIA VIAG1_N_WW
  LAYER MET5 ;
    RECT -0.260 -0.200 0.260 0.320 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.140 0.200 0.260 ;
  LAYER METG1 ;
    RECT -0.200 -0.140 0.200 0.260 ;
END VIAG1_N_WW

VIA VIAG1_S_WW
  LAYER MET5 ;
    RECT -0.260 -0.320 0.260 0.200 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.260 0.200 0.140 ;
  LAYER METG1 ;
    RECT -0.200 -0.260 0.200 0.140 ;
END VIAG1_S_WW

VIA VIAG1_E_WW
  LAYER MET5 ;
    RECT -0.200 -0.260 0.320 0.260 ;
  LAYER CUTG1 ;
    RECT -0.140 -0.200 0.260 0.200 ;
  LAYER METG1 ;
    RECT -0.140 -0.200 0.260 0.200 ;
END VIAG1_E_WW

VIA VIAG1_W_WW
  LAYER MET5 ;
    RECT -0.320 -0.260 0.200 0.260 ;
  LAYER CUTG1 ;
    RECT -0.260 -0.200 0.140 0.200 ;
  LAYER METG1 ;
    RECT -0.260 -0.200 0.140 0.200 ;
END VIAG1_W_WW

# MULTI-VIA
VIA VIAG1_2N_WW
  LAYER MET5 ;
    RECT -0.260 -0.260 0.260 1.060 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
    RECT -0.200  0.600 0.200 1.000 ;
  LAYER METG1 ;
    RECT -0.200 -0.200 0.200 1.000 ;
END VIAG1_2N_WW

VIA VIAG1_2S_WW
  LAYER MET5 ;
    RECT -0.260 -1.060 0.260  0.260 ;
  LAYER CUTG1 ;
    RECT -0.200 -1.000 0.200 -0.600 ;
    RECT -0.200 -0.200 0.200  0.200 ;
  LAYER METG1 ;
    RECT -0.200 -1.000 0.200  0.200 ;
END VIAG1_2S_WW

VIA VIAG1_2V_WW
  LAYER MET5 ;
    RECT -0.260 -0.660 0.260  0.660 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.600 0.200 -0.200 ;
    RECT -0.200  0.200 0.200  0.600 ;
  LAYER METG1 ;
    RECT -0.200 -0.600 0.200  0.600 ;
END VIAG1_2V_WW

VIA VIAG1_2E_WW
  LAYER MET5 ;
    RECT -0.260 -0.260 1.060  0.260 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200  0.200 ;
    RECT  0.600 -0.200 1.000  0.200 ;
  LAYER METG1 ;
    RECT -0.200 -0.200 1.000  0.200 ;
END VIAG1_2E_WW

VIA VIAG1_2W_WW
  LAYER MET5 ;
    RECT -1.060 -0.260  0.260 0.260 ;
  LAYER CUTG1 ;
    RECT -1.000 -0.200 -0.600 0.200 ;
    RECT -0.200 -0.200  0.200 0.200 ;
  LAYER METG1 ;
    RECT -1.000 -0.200  0.200 0.200 ;
END VIAG1_2W_WW

VIA VIAG1_2H_WW
  LAYER MET5 ;
    RECT -0.660 -0.260  0.660 0.260 ;
  LAYER CUTG1 ;
    RECT -0.600 -0.200 -0.200 0.200 ;
    RECT  0.200 -0.200  0.600 0.200 ;
  LAYER METG1 ;
    RECT -0.600 -0.200  0.600 0.200 ;
END VIAG1_2H_WW

# SINGLE/STACK-VIA
VIA VIATOP_WW
  LAYER METG1 ;
    RECT -0.350 -0.350 0.350 0.350 ;
  LAYER CUTTOP ;
    RECT -0.250 -0.250 0.250 0.250 ;
  LAYER METTOP ;
    RECT -0.500 -0.500 0.500 0.500 ;
END VIATOP_WW

# MULTI-VIA
VIA VIATOP_2N_WW
  LAYER METG1 ;
    RECT -0.350 -0.350 0.350 1.950 ;
  LAYER CUTTOP ;
    RECT -0.250 -0.250 0.250 0.250 ;
    RECT -0.250  1.350 0.250 1.850 ;
  LAYER METTOP ;
    RECT -0.500 -0.500 0.500 2.100 ;
END VIATOP_2N_WW

VIA VIATOP_2S_WW
  LAYER METG1 ;
    RECT -0.350 -1.950 0.350  0.350 ;
  LAYER CUTTOP ;
    RECT -0.250 -1.850 0.250 -1.350 ;
    RECT -0.250 -0.250 0.250  0.250 ;
  LAYER METTOP ;
    RECT -0.500 -2.100 0.500  0.500 ;
END VIATOP_2S_WW

VIA VIATOP_2V_WW
  LAYER METG1 ;
    RECT -0.350 -1.150 0.350  1.150 ;
  LAYER CUTTOP ;
    RECT -0.250 -1.050 0.250 -0.550 ;
    RECT -0.250  0.550 0.250  1.050 ;
  LAYER METTOP ;
    RECT -0.500 -1.300 0.500  1.300 ;
END VIATOP_2V_WW

VIA VIATOP_2E_WW
  LAYER METG1 ;
    RECT -0.350 -0.350 1.950 0.350 ;
  LAYER CUTTOP ;
    RECT -0.250 -0.250 0.250 0.250 ;
    RECT  1.350 -0.250 1.850 0.250 ;
  LAYER METTOP ;
    RECT -0.500 -0.500 2.100 0.500 ;
END VIATOP_2E_WW

VIA VIATOP_2W_WW
  LAYER METG1 ;
    RECT -1.950 -0.350  0.350 0.350 ;
  LAYER CUTTOP ;
    RECT -1.850 -0.250 -1.350 0.250 ;
    RECT -0.250 -0.250  0.250 0.250 ;
  LAYER METTOP ;
    RECT -2.100 -0.500  0.500 0.500 ;
END VIATOP_2W_WW

VIA VIATOP_2H_WW
  LAYER METG1 ;
    RECT -1.150 -0.350  1.150 0.350 ;
  LAYER CUTTOP ;
    RECT -1.050 -0.250 -0.550 0.250 ;
    RECT  0.550 -0.250  1.050 0.250 ;
  LAYER METTOP ;
    RECT -1.300 -0.500  1.300 0.500 ;
END VIATOP_2H_WW

END WIDEWIRE

NONDEFAULTRULE WIDEWIRE_DC
LAYER MET1
  WIDTH 0.100 ;
  SPACING 0.100 ;
END MET1

LAYER MET2
  WIDTH 0.100 ;
  SPACING 0.100 ;
END MET2

LAYER MET3
  WIDTH 0.100 ;
  SPACING 0.100 ;
END MET3

LAYER MET4
  WIDTH 0.180 ;
  SPACING 0.120 ;
END MET4

LAYER MET5
  WIDTH 0.180 ;
  SPACING 0.120 ;
END MET5

LAYER METG1
  WIDTH 0.400 ;
  SPACING 0.400 ;
END METG1

LAYER METTOP
  WIDTH 0.800 ;
  SPACING 0.800 ;
END METTOP

# MULTI-VIA
VIA VIA1_2N_WWDC
  LAYER MET1 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA1_2N_WWDC

VIA VIA1_2NV_WWDC
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA1_2NV_WWDC

VIA VIA1_2NR_WWDC
  LAYER MET1 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA1_2NR_WWDC

VIA VIA1_2S_WWDC
  LAYER MET1 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA1_2S_WWDC

VIA VIA1_2SV_WWDC
  LAYER MET1 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA1_2SV_WWDC

VIA VIA1_2SR_WWDC
  LAYER MET1 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA1_2SR_WWDC

VIA VIA1_2V_WWDC
  LAYER MET1 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA1_2V_WWDC

VIA VIA1_2CV_WWDC
  LAYER MET1 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA1_2CV_WWDC

VIA VIA1_2VR_WWDC
  LAYER MET1 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT12 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET2 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA1_2VR_WWDC

VIA VIA1_2E_WWDC
  LAYER MET1 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA1_2E_WWDC

VIA VIA1_2EH_WWDC
  LAYER MET1 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA1_2EH_WWDC

VIA VIA1_2ER_WWDC
  LAYER MET1 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA1_2ER_WWDC

VIA VIA1_2W_WWDC
  LAYER MET1 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA1_2W_WWDC

VIA VIA1_2WH_WWDC
  LAYER MET1 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA1_2WH_WWDC

VIA VIA1_2WR_WWDC
  LAYER MET1 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA1_2WR_WWDC

VIA VIA1_2H_WWDC
  LAYER MET1 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA1_2H_WWDC

VIA VIA1_2CH_WWDC
  LAYER MET1 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA1_2CH_WWDC

VIA VIA1_2HR_WWDC
  LAYER MET1 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT12 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA1_2HR_WWDC

VIA VIA1_3H_WWDC
  LAYER MET1 ;
    RECT -0.290 -0.050  0.290 0.050 ;
  LAYER CUT12 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET2 ;
    RECT -0.250 -0.090  0.250 0.090 ;
END VIA1_3H_WWDC

VIA VIA1_3V_WWDC
  LAYER MET1 ;
    RECT -0.090 -0.250 0.090  0.250 ;
  LAYER CUT12 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.290 ;
END VIA1_3V_WWDC

VIA VIA1_4H_WWDC
  LAYER MET1 ;
    RECT -0.390 -0.050  0.390 0.050 ;
  LAYER CUT12 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET2 ;
    RECT -0.350 -0.090  0.350 0.090 ;
END VIA1_4H_WWDC

VIA VIA1_4V_WWDC
  LAYER MET1 ;
    RECT -0.090 -0.350 0.090  0.350 ;
  LAYER CUT12 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET2 ;
    RECT -0.050 -0.390 0.050  0.390 ;
END VIA1_4V_WWDC

# MULTI-VIA
VIA VIA2_2N_WWDC
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA2_2N_WWDC

VIA VIA2_2NV_WWDC
  LAYER MET2 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA2_2NV_WWDC

VIA VIA2_2NR_WWDC
  LAYER MET2 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
END VIA2_2NR_WWDC

VIA VIA2_2S_WWDC
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA2_2S_WWDC

VIA VIA2_2SV_WWDC
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA2_2SV_WWDC

VIA VIA2_2SR_WWDC
  LAYER MET2 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
END VIA2_2SR_WWDC

VIA VIA2_2V_WWDC
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA2_2V_WWDC

VIA VIA2_2CV_WWDC
  LAYER MET2 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA2_2CV_WWDC

VIA VIA2_2VR_WWDC
  LAYER MET2 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT23 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
END VIA2_2VR_WWDC

VIA VIA2_2E_WWDC
  LAYER MET2 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA2_2E_WWDC

VIA VIA2_2EH_WWDC
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
END VIA2_2EH_WWDC

VIA VIA2_2ER_WWDC
  LAYER MET2 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA2_2ER_WWDC

VIA VIA2_2W_WWDC
  LAYER MET2 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA2_2W_WWDC

VIA VIA2_2WH_WWDC
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
END VIA2_2WH_WWDC

VIA VIA2_2WR_WWDC
  LAYER MET2 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET3 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA2_2WR_WWDC

VIA VIA2_2H_WWDC
  LAYER MET2 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA2_2H_WWDC

VIA VIA2_2CH_WWDC
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.190 -0.050  0.190 0.050 ;
END VIA2_2CH_WWDC

VIA VIA2_2HR_WWDC
  LAYER MET2 ;
    RECT -0.190 -0.050  0.190 0.050 ;
  LAYER CUT23 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET3 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA2_2HR_WWDC

VIA VIA2_3H_WWDC
  LAYER MET2 ;
    RECT -0.250 -0.090  0.250 0.090 ;
  LAYER CUT23 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET3 ;
    RECT -0.290 -0.050  0.290 0.050 ;
END VIA2_3H_WWDC

VIA VIA2_3V_WWDC
  LAYER MET2 ;
    RECT -0.050 -0.290 0.050  0.290 ;
  LAYER CUT23 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.250 ;
END VIA2_3V_WWDC

VIA VIA2_4H_WWDC
  LAYER MET2 ;
    RECT -0.350 -0.090  0.350 0.090 ;
  LAYER CUT23 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET3 ;
    RECT -0.390 -0.050  0.390 0.050 ;
END VIA2_4H_WWDC

VIA VIA2_4V_WWDC
  LAYER MET2 ;
    RECT -0.050 -0.390 0.050  0.390 ;
  LAYER CUT23 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET3 ;
    RECT -0.090 -0.350 0.090  0.350 ;
END VIA2_4V_WWDC

# MULTI-VIA
VIA VIA3_2N_WWDC
  LAYER MET3 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA3_2N_WWDC

VIA VIA3_2S_WWDC
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA3_2S_WWDC

VIA VIA3_2E_WWDC
  LAYER MET3 ;
    RECT -0.090 -0.050 0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA3_2E_WWDC

VIA VIA3_2W_WWDC
  LAYER MET3 ;
    RECT -0.290 -0.050  0.090 0.050 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA3_2W_WWDC

VIA VIA3_2NR_WWDC
  LAYER MET3 ;
    RECT -0.050 -0.090 0.050 0.290 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA3_2NR_WWDC

VIA VIA3_2SR_WWDC
  LAYER MET3 ;
    RECT -0.050 -0.290 0.050  0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA3_2SR_WWDC

VIA VIA3_2ER_WWDC
  LAYER MET3 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA3_2ER_WWDC

VIA VIA3_2WR_WWDC
  LAYER MET3 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET4 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA3_2WR_WWDC

VIA VIA3_2CH_WWDC
  LAYER MET3 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT34 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET4 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA3_2CH_WWDC

VIA VIA3_2VR_WWDC
  LAYER MET3 ;
    RECT -0.050 -0.190 0.050  0.190 ;
  LAYER CUT34 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET4 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA3_2VR_WWDC

VIA VIA3_3H_WWDC
  LAYER MET3 ;
    RECT -0.290 -0.050  0.290 0.050 ;
  LAYER CUT34 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET4 ;
    RECT -0.250 -0.090  0.250 0.090 ;
END VIA3_3H_WWDC

VIA VIA3_3V_WWDC
  LAYER MET3 ;
    RECT -0.090 -0.250 0.090  0.250 ;
  LAYER CUT34 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.250 ;
END VIA3_3V_WWDC

VIA VIA3_4H_WWDC
  LAYER MET3 ;
    RECT -0.390 -0.050  0.390 0.050 ;
  LAYER CUT34 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET4 ;
    RECT -0.350 -0.090  0.350 0.090 ;
END VIA3_4H_WWDC

VIA VIA3_4V_WWDC
  LAYER MET3 ;
    RECT -0.090 -0.350 0.090  0.350 ;
  LAYER CUT34 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET4 ;
    RECT -0.090 -0.350 0.090  0.350 ;
END VIA3_4V_WWDC

# MULTI-VIA
VIA VIA4_2N_WWDC
  LAYER MET4 ;
    RECT -0.090 -0.050 0.090 0.250 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT -0.050  0.150 0.050 0.250 ;
  LAYER MET5 ;
    RECT -0.090 -0.050 0.090 0.250 ;
END VIA4_2N_WWDC

VIA VIA4_2S_WWDC
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.050 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
  LAYER MET5 ;
    RECT -0.090 -0.250 0.090  0.050 ;
END VIA4_2S_WWDC

VIA VIA4_2V_WWDC
  LAYER MET4 ;
    RECT -0.090 -0.150 0.090  0.150 ;
  LAYER CUT45 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
  LAYER MET5 ;
    RECT -0.090 -0.150 0.090  0.150 ;
END VIA4_2V_WWDC

VIA VIA4_2E_WWDC
  LAYER MET4 ;
    RECT -0.050 -0.090 0.250 0.090 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    RECT  0.150 -0.050 0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.050 -0.090 0.250 0.090 ;
END VIA4_2E_WWDC

VIA VIA4_2W_WWDC
  LAYER MET4 ;
    RECT -0.250 -0.090  0.050 0.090 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
  LAYER MET5 ;
    RECT -0.250 -0.090  0.050 0.090 ;
END VIA4_2W_WWDC

VIA VIA4_2H_WWDC
  LAYER MET4 ;
    RECT -0.150 -0.090  0.150 0.090 ;
  LAYER CUT45 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
  LAYER MET5 ;
    RECT -0.150 -0.090  0.150 0.090 ;
END VIA4_2H_WWDC

VIA VIA4_3H_WWDC
  LAYER MET4 ;
    RECT -0.250 -0.090  0.250 0.090 ;
  LAYER CUT45 ;
    RECT -0.250 -0.050 -0.150 0.050 ;
    RECT -0.050 -0.050  0.050 0.050 ;
    RECT  0.150 -0.050  0.250 0.050 ;
  LAYER MET5 ;
    RECT -0.250 -0.090  0.250 0.090 ;
END VIA4_3H_WWDC

VIA VIA4_3V_WWDC
  LAYER MET4 ;
    RECT -0.090 -0.250 0.090  0.250 ;
  LAYER CUT45 ;
    RECT -0.050 -0.250 0.050 -0.150 ;
    RECT -0.050 -0.050 0.050  0.050 ;
    RECT -0.050  0.150 0.050  0.250 ;
  LAYER MET5 ;
    RECT -0.090 -0.250 0.090  0.250 ;
END VIA4_3V_WWDC

VIA VIA4_4H_WWDC
  LAYER MET4 ;
    RECT -0.350 -0.090  0.350 0.090 ;
  LAYER CUT45 ;
    RECT -0.350 -0.050 -0.250 0.050 ;
    RECT -0.150 -0.050 -0.050 0.050 ;
    RECT  0.050 -0.050  0.150 0.050 ;
    RECT  0.250 -0.050  0.350 0.050 ;
  LAYER MET5 ;
    RECT -0.350 -0.090  0.350 0.090 ;
END VIA4_4H_WWDC

VIA VIA4_4V_WWDC
  LAYER MET4 ;
    RECT -0.090 -0.350 0.090  0.350 ;
  LAYER CUT45 ;
    RECT -0.050 -0.350 0.050 -0.250 ;
    RECT -0.050 -0.150 0.050 -0.050 ;
    RECT -0.050  0.050 0.050  0.150 ;
    RECT -0.050  0.250 0.050  0.350 ;
  LAYER MET5 ;
    RECT -0.090 -0.350 0.090  0.350 ;
END VIA4_4V_WWDC

# MULTI-VIA
VIA VIAG1_2N_WWDC
  LAYER MET5 ;
    RECT -0.260 -0.260 0.260 1.060 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
    RECT -0.200  0.600 0.200 1.000 ;
  LAYER METG1 ;
    RECT -0.200 -0.200 0.200 1.000 ;
END VIAG1_2N_WWDC

VIA VIAG1_2S_WWDC
  LAYER MET5 ;
    RECT -0.260 -1.060 0.260  0.260 ;
  LAYER CUTG1 ;
    RECT -0.200 -1.000 0.200 -0.600 ;
    RECT -0.200 -0.200 0.200  0.200 ;
  LAYER METG1 ;
    RECT -0.200 -1.000 0.200  0.200 ;
END VIAG1_2S_WWDC

VIA VIAG1_2V_WWDC
  LAYER MET5 ;
    RECT -0.260 -0.660 0.260  0.660 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.600 0.200 -0.200 ;
    RECT -0.200  0.200 0.200  0.600 ;
  LAYER METG1 ;
    RECT -0.200 -0.600 0.200  0.600 ;
END VIAG1_2V_WWDC

VIA VIAG1_2E_WWDC
  LAYER MET5 ;
    RECT -0.260 -0.260 1.060  0.260 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200  0.200 ;
    RECT  0.600 -0.200 1.000  0.200 ;
  LAYER METG1 ;
    RECT -0.200 -0.200 1.000  0.200 ;
END VIAG1_2E_WWDC

VIA VIAG1_2W_WWDC
  LAYER MET5 ;
    RECT -1.060 -0.260  0.260 0.260 ;
  LAYER CUTG1 ;
    RECT -1.000 -0.200 -0.600 0.200 ;
    RECT -0.200 -0.200  0.200 0.200 ;
  LAYER METG1 ;
    RECT -1.000 -0.200  0.200 0.200 ;
END VIAG1_2W_WWDC

VIA VIAG1_2H_WWDC
  LAYER MET5 ;
    RECT -0.660 -0.260  0.660 0.260 ;
  LAYER CUTG1 ;
    RECT -0.600 -0.200 -0.200 0.200 ;
    RECT  0.200 -0.200  0.600 0.200 ;
  LAYER METG1 ;
    RECT -0.600 -0.200  0.600 0.200 ;
END VIAG1_2H_WWDC

# MULTI-VIA
VIA VIATOP_2N_WWDC
  LAYER METG1 ;
    RECT -0.350 -0.350 0.350 1.950 ;
  LAYER CUTTOP ;
    RECT -0.250 -0.250 0.250 0.250 ;
    RECT -0.250  1.350 0.250 1.850 ;
  LAYER METTOP ;
    RECT -0.500 -0.500 0.500 2.100 ;
END VIATOP_2N_WWDC

VIA VIATOP_2S_WWDC
  LAYER METG1 ;
    RECT -0.350 -1.950 0.350  0.350 ;
  LAYER CUTTOP ;
    RECT -0.250 -1.850 0.250 -1.350 ;
    RECT -0.250 -0.250 0.250  0.250 ;
  LAYER METTOP ;
    RECT -0.500 -2.100 0.500  0.500 ;
END VIATOP_2S_WWDC

VIA VIATOP_2V_WWDC
  LAYER METG1 ;
    RECT -0.350 -1.150 0.350  1.150 ;
  LAYER CUTTOP ;
    RECT -0.250 -1.050 0.250 -0.550 ;
    RECT -0.250  0.550 0.250  1.050 ;
  LAYER METTOP ;
    RECT -0.500 -1.300 0.500  1.300 ;
END VIATOP_2V_WWDC

VIA VIATOP_2E_WWDC
  LAYER METG1 ;
    RECT -0.350 -0.350 1.950 0.350 ;
  LAYER CUTTOP ;
    RECT -0.250 -0.250 0.250 0.250 ;
    RECT  1.350 -0.250 1.850 0.250 ;
  LAYER METTOP ;
    RECT -0.500 -0.500 2.100 0.500 ;
END VIATOP_2E_WWDC

VIA VIATOP_2W_WWDC
  LAYER METG1 ;
    RECT -1.950 -0.350  0.350 0.350 ;
  LAYER CUTTOP ;
    RECT -1.850 -0.250 -1.350 0.250 ;
    RECT -0.250 -0.250  0.250 0.250 ;
  LAYER METTOP ;
    RECT -2.100 -0.500  0.500 0.500 ;
END VIATOP_2W_WWDC

VIA VIATOP_2H_WWDC
  LAYER METG1 ;
    RECT -1.150 -0.350  1.150 0.350 ;
  LAYER CUTTOP ;
    RECT -1.050 -0.250 -0.550 0.250 ;
    RECT  0.550 -0.250  1.050 0.250 ;
  LAYER METTOP ;
    RECT -1.300 -0.500  1.300 0.500 ;
END VIATOP_2H_WWDC

END WIDEWIRE_DC

# === LEF v5.5 SPEC ===
#VIARULE TURNMET1 GENERATE
#  LAYER MET1 ;
#    DIRECTION VERTICAL ;
#  LAYER MET1 ;
#    DIRECTION HORIZONTAL ;
#END TURNMET1
# === END ===

# === LEF v5.5 SPEC ===
#VIARULE TURNMET2 GENERATE
#  LAYER MET2 ;
#    DIRECTION VERTICAL ;
#  LAYER MET2 ;
#    DIRECTION HORIZONTAL ;
#END TURNMET2
# === END ===

# === LEF v5.5 SPEC ===
#VIARULE TURNMET3 GENERATE
#  LAYER MET3 ;
#    DIRECTION VERTICAL ;
#  LAYER MET3 ;
#    DIRECTION HORIZONTAL ;
#END TURNMET3
# === END ===

# === LEF v5.5 SPEC ===
#VIARULE TURNMET4 GENERATE
#  LAYER MET4 ;
#    DIRECTION VERTICAL ;
#  LAYER MET4 ;
#    DIRECTION HORIZONTAL ;
#END TURNMET4
# === END ===

# === LEF v5.5 SPEC ===
#VIARULE TURNMET5 GENERATE
#  LAYER MET5 ;
#    DIRECTION VERTICAL ;
#  LAYER MET5 ;
#    DIRECTION HORIZONTAL ;
#END TURNMET5
# === END ===

# === LEF v5.5 SPEC ===
#VIARULE TURNMETG1 GENERATE
#  LAYER METG1 ;
#    DIRECTION VERTICAL ;
#  LAYER METG1 ;
#    DIRECTION HORIZONTAL ;
#END TURNMETG1
# === END ===

# === LEF v5.5 SPEC ===
#VIARULE TURNMETTOP GENERATE
#  LAYER METTOP ;
#    DIRECTION VERTICAL ;
#  LAYER METTOP ;
#    DIRECTION HORIZONTAL ;
#END TURNMETTOP
# === END ===

VIARULE VIAGEN11 GENERATE
  LAYER MET1 ;
    WIDTH 0.100 TO 0.500 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER MET2 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN11

VIARULE VIAGEN12 GENERATE
  LAYER MET1 ;
    WIDTH 0.100 TO 0.500 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER MET2 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN12

VIARULE VIAGEN13 GENERATE
  LAYER MET1 ;
    WIDTH 0.100 TO 0.500 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER MET2 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN13

VIARULE VIAGEN14 GENERATE
  LAYER MET1 ;
    WIDTH 0.501 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER MET2 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN14

VIARULE VIAGEN15 GENERATE
  LAYER MET1 ;
    WIDTH 0.501 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER MET2 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN15

VIARULE VIAGEN16 GENERATE
  LAYER MET1 ;
    WIDTH 0.501 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER MET2 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN16

VIARULE VIAGEN17 GENERATE
  LAYER MET1 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER MET2 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN17

VIARULE VIAGEN18 GENERATE
  LAYER MET1 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER MET2 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN18

VIARULE VIAGEN19 GENERATE
  LAYER MET1 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER MET2 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER CUT12 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN19

VIARULE VIAGEN21 GENERATE
  LAYER MET2 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER MET3 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN21

VIARULE VIAGEN22 GENERATE
  LAYER MET2 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER MET3 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN22

VIARULE VIAGEN23 GENERATE
  LAYER MET2 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER MET3 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN23

VIARULE VIAGEN24 GENERATE
  LAYER MET2 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER MET3 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN24

VIARULE VIAGEN25 GENERATE
  LAYER MET2 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER MET3 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN25

VIARULE VIAGEN26 GENERATE
  LAYER MET2 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER MET3 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN26

VIARULE VIAGEN27 GENERATE
  LAYER MET2 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER MET3 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN27

VIARULE VIAGEN28 GENERATE
  LAYER MET2 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER MET3 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN28

VIARULE VIAGEN29 GENERATE
  LAYER MET2 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER MET3 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER CUT23 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN29

# POWER-RAIL VIA
VIARULE VIARULE341
  LAYER MET3 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.300 TO 0.300 ;
  LAYER MET4 ;
    DIRECTION VERTICAL ;
    WIDTH 1.450 TO 1.450 ;
  VIA VIA34P ;
END VIARULE341

# POWER-RAIL VIA
VIARULE VIARULE342
  LAYER MET3 ;
    DIRECTION HORIZONTAL ;
    WIDTH 0.320 TO 0.320 ;
  LAYER MET4 ;
    DIRECTION VERTICAL ;
    WIDTH 1.450 TO 1.450 ;
  VIA VIA34P2 ;
END VIARULE342

VIARULE VIAGEN31 GENERATE
  LAYER MET3 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER MET4 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN31

VIARULE VIAGEN32 GENERATE
  LAYER MET3 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER MET4 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN32

VIARULE VIAGEN33 GENERATE
  LAYER MET3 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER MET4 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN33

VIARULE VIAGEN34 GENERATE
  LAYER MET3 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER MET4 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN34

VIARULE VIAGEN35 GENERATE
  LAYER MET3 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER MET4 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN35

VIARULE VIAGEN36 GENERATE
  LAYER MET3 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER MET4 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN36

VIARULE VIAGEN37 GENERATE
  LAYER MET3 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER MET4 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN37

VIARULE VIAGEN38 GENERATE
  LAYER MET3 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER MET4 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN38

VIARULE VIAGEN39 GENERATE
  LAYER MET3 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER MET4 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER CUT34 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN39

VIARULE VIAGEN41 GENERATE
  LAYER MET4 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER MET5 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN41

VIARULE VIAGEN42 GENERATE
  LAYER MET4 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER MET5 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN42

VIARULE VIAGEN43 GENERATE
  LAYER MET4 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER MET5 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN43

VIARULE VIAGEN44 GENERATE
  LAYER MET4 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER MET5 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN44

VIARULE VIAGEN45 GENERATE
  LAYER MET4 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER MET5 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN45

VIARULE VIAGEN46 GENERATE
  LAYER MET4 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER MET5 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN46

VIARULE VIAGEN47 GENERATE
  LAYER MET4 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER MET5 ;
    WIDTH 0.100 TO 0.800 ;
    ENCLOSURE 0.000 0.040 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN47

VIARULE VIAGEN48 GENERATE
  LAYER MET4 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER MET5 ;
    WIDTH 0.801 TO 1.200 ;
    ENCLOSURE 0.015 0.040 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN48

VIARULE VIAGEN49 GENERATE
  LAYER MET4 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER MET5 ;
    WIDTH 1.201 TO 1000.000 ;
    ENCLOSURE 0.035 0.040 ;
  LAYER CUT45 ;
    RECT -0.050 -0.050 0.050 0.050 ;
    SPACING 0.200 by 0.200 ;
END VIAGEN49

VIARULE VIAGENG11 GENERATE
  LAYER MET5 ;
    WIDTH 0.100 TO 1.260 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER METG1 ;
    WIDTH 0.400 TO 1.400 ;
    ENCLOSURE 0.000 0.000 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
    SPACING 0.800 by 0.800 ;
END VIAGENG11

VIARULE VIAGENG12 GENERATE
  LAYER MET5 ;
    WIDTH 0.100 TO 1.260 ;
    ENCLOSURE 0.060 0.060 ;
  LAYER METG1 ;
    WIDTH 1.401 TO 1000.000 ;
    ENCLOSURE 0.100 0.100 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
    SPACING 0.800 by 0.800 ;
END VIAGENG12

VIARULE VIAGENG13 GENERATE
  LAYER MET5 ;
    WIDTH 1.261 TO 1000.000 ;
    ENCLOSURE 0.100 0.100 ;
  LAYER METG1 ;
    WIDTH 0.400 TO 1.400 ;
    ENCLOSURE 0.000 0.000 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
    SPACING 0.800 by 0.800 ;
END VIAGENG13

VIARULE VIAGENG14 GENERATE
  LAYER MET5 ;
    WIDTH 1.261 TO 1000.000 ;
    ENCLOSURE 0.100 0.100 ;
  LAYER METG1 ;
    WIDTH 1.401 TO 1000.000 ;
    ENCLOSURE 0.100 0.100 ;
  LAYER CUTG1 ;
    RECT -0.200 -0.200 0.200 0.200 ;
    SPACING 0.800 by 0.800 ;
END VIAGENG14

VIARULE VIAGENTOP GENERATE
  LAYER METG1 ;
    WIDTH 0.400 TO 1000.000 ;
    ENCLOSURE 0.100 0.100 ;
  LAYER METTOP ;
    WIDTH 0.800 TO 1000.000 ;
    ENCLOSURE 0.250 0.250 ;
  LAYER CUTTOP ;
    RECT -0.250 -0.250 0.250 0.250 ;
    SPACING 1.600 by 1.600 ;
END VIAGENTOP

SITE COVER
  CLASS PAD ;
  SIZE 1 BY 1 ;
END COVER

END LIBRARY